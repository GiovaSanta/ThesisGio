--------------------------------------------------------------------------------
--                            MultTable_comb_uid7_fixP16_32 # i renamed it because the old name was used also in the 
--                                          fixed point 8_16  MAC module
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid7_fixP16_32 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid7_fixP16_32 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "010" when "101",
      "000" when "110",
      "001" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid11
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid11 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid11 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "11110" when "10001",
      "11100" when "10010",
      "11010" when "10011",
      "11000" when "10100",
      "10110" when "10101",
      "10100" when "10110",
      "10010" when "10111",
      "00000" when "11000",
      "11111" when "11001",
      "11110" when "11010",
      "11101" when "11011",
      "11100" when "11100",
      "11011" when "11101",
      "11010" when "11110",
      "11001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid15
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid15 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid15 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "11110" when "10001",
      "11100" when "10010",
      "11010" when "10011",
      "11000" when "10100",
      "10110" when "10101",
      "10100" when "10110",
      "10010" when "10111",
      "00000" when "11000",
      "11111" when "11001",
      "11110" when "11010",
      "11101" when "11011",
      "11100" when "11100",
      "11011" when "11101",
      "11010" when "11110",
      "11001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid19
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid19 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid19 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "11110" when "10001",
      "11100" when "10010",
      "11010" when "10011",
      "11000" when "10100",
      "10110" when "10101",
      "10100" when "10110",
      "10010" when "10111",
      "00000" when "11000",
      "11111" when "11001",
      "11110" when "11010",
      "11101" when "11011",
      "11100" when "11100",
      "11011" when "11101",
      "11010" when "11110",
      "11001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid23
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid23 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid23 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "11110" when "10001",
      "11100" when "10010",
      "11010" when "10011",
      "11000" when "10100",
      "10110" when "10101",
      "10100" when "10110",
      "10010" when "10111",
      "00000" when "11000",
      "11111" when "11001",
      "11110" when "11010",
      "11101" when "11011",
      "11100" when "11100",
      "11011" when "11101",
      "11010" when "11110",
      "11001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid27
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "11110" when "10001",
      "11100" when "10010",
      "11010" when "10011",
      "11000" when "10100",
      "10110" when "10101",
      "10100" when "10110",
      "10010" when "10111",
      "00000" when "11000",
      "11111" when "11001",
      "11110" when "11010",
      "11101" when "11011",
      "11100" when "11100",
      "11011" when "11101",
      "11010" when "11110",
      "11001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid31
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid31 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid31 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid35
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid35 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid35 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid39
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid39 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid39 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid43
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid43 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid43 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid47
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid47 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid47 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid51
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid51 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid51 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid55
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid55 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid55 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid59
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid59 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid59 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid63
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid67
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid67 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid67 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid71
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid71 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid71 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid75
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid75 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid75 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid79
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid79 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid79 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid83
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid87
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid87 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid87 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid91
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid91 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid91 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid95
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid95 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid95 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_comb_uid99
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid99 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid99 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid103
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid103 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid103 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid107
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid107 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid107 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid111
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid111 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid111 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid115
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid115 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid115 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid119
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid119 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid119 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid123
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid127
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid127 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid127 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid131
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid131 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid131 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid135
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid135 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid135 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid139
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid139 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid139 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid143
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid143 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid143 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid147
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid147 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid147 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid151
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid151 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid151 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid155
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid155 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid155 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid159
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid159 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid159 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid163
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid163 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid163 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid167
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid167 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid167 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid171
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid171 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid171 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid175
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid175 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid175 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000",
      "000" when "001",
      "000" when "010",
      "111" when "011",
      "000" when "100",
      "110" when "101",
      "000" when "110",
      "101" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid179
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid179 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid179 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid183
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid183 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid183 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid187
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid187 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid187 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid191
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid191 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid191 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_comb_uid195
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_comb_uid195 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_comb_uid195 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_23_3_comb_uid198
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_comb_uid198 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_comb_uid198 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_3_2_comb_uid201
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_comb_uid201 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_comb_uid201 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_14_3_comb_uid204
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_comb_uid204 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_comb_uid204 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_6_3_comb_uid209
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_comb_uid209 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_comb_uid209 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_1_signedx2_signed_comb_uid5
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_signed_comb_uid5 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_signed_comb_uid5 is
   component MultTable_comb_uid7_fixP16_32 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid7_fixP16_32
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_3x2_signed_comb_uid9
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_signed_comb_uid9 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_signed_comb_uid9 is
   component MultTable_comb_uid11 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid11
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_3x2_signed_comb_uid13
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_signed_comb_uid13 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_signed_comb_uid13 is
   component MultTable_comb_uid15 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid15
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_3x2_signed_comb_uid17
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_signed_comb_uid17 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_signed_comb_uid17 is
   component MultTable_comb_uid19 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid19
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_3x2_signed_comb_uid21
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_signed_comb_uid21 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_signed_comb_uid21 is
   component MultTable_comb_uid23 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid23
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_3x2_signed_comb_uid25
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_signed_comb_uid25 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_signed_comb_uid25 is
   component MultTable_comb_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid27
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_1_signedx2_comb_uid29
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid29 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid29 is
   component MultTable_comb_uid31 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid31
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid33
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid33 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid33 is
   component MultTable_comb_uid35 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid35
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid37
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid37 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid37 is
   component MultTable_comb_uid39 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid39
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid41
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid41 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid41 is
   component MultTable_comb_uid43 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid43
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid45
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid45 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid45 is
   component MultTable_comb_uid47 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid47
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid49
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid49 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid49 is
   component MultTable_comb_uid51 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid51
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_1_signedx2_comb_uid53
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid53 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid53 is
   component MultTable_comb_uid55 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid55
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid57
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid57 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid57 is
   component MultTable_comb_uid59 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid59
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid61
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid61 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid61 is
   component MultTable_comb_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid63
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid65
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid65 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid65 is
   component MultTable_comb_uid67 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid67
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid69
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid69 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid69 is
   component MultTable_comb_uid71 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid71
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid73
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid73 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid73 is
   component MultTable_comb_uid75 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid75
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplierLUT_1_signedx2_comb_uid77
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid77 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid77 is
   component MultTable_comb_uid79 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid79
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid81
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid81 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid81 is
   component MultTable_comb_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid83
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid85
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid85 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid85 is
   component MultTable_comb_uid87 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid87
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid89
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid89 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid89 is
   component MultTable_comb_uid91 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid91
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid93
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid93 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid93 is
   component MultTable_comb_uid95 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid95
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid97
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid97 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid97 is
   component MultTable_comb_uid99 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid99
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                  IntMultiplierLUT_1_signedx2_comb_uid101
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid101 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid101 is
   component MultTable_comb_uid103 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid103
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid105
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid105 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid105 is
   component MultTable_comb_uid107 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid107
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid109
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid109 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid109 is
   component MultTable_comb_uid111 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid111
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid113
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid113 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid113 is
   component MultTable_comb_uid115 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid115
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid117
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid117 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid117 is
   component MultTable_comb_uid119 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid119
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid121
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid121 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid121 is
   component MultTable_comb_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid123
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                  IntMultiplierLUT_1_signedx2_comb_uid125
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid125 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid125 is
   component MultTable_comb_uid127 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid127
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid129
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid129 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid129 is
   component MultTable_comb_uid131 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid131
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid133
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid133 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid133 is
   component MultTable_comb_uid135 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid135
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid137
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid137 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid137 is
   component MultTable_comb_uid139 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid139
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid141
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid141 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid141 is
   component MultTable_comb_uid143 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid143
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid145
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid145 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid145 is
   component MultTable_comb_uid147 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid147
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                  IntMultiplierLUT_1_signedx2_comb_uid149
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid149 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid149 is
   component MultTable_comb_uid151 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid151
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid153
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid153 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid153 is
   component MultTable_comb_uid155 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid155
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid157
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid157 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid157 is
   component MultTable_comb_uid159 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid159
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid161
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid161 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid161 is
   component MultTable_comb_uid163 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid163
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid165
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid165 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid165 is
   component MultTable_comb_uid167 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid167
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid169
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid169 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid169 is
   component MultTable_comb_uid171 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid171
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                  IntMultiplierLUT_1_signedx2_comb_uid173
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1_signedx2_comb_uid173 is
    port (X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1_signedx2_comb_uid173 is
   component MultTable_comb_uid175 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(2 downto 0);
signal Y1 :  std_logic_vector(2 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid175
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid177
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid177 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid177 is
   component MultTable_comb_uid179 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid179
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid181
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid181 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid181 is
   component MultTable_comb_uid183 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid183
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid185
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid185 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid185 is
   component MultTable_comb_uid187 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid187
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid189
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid189 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid189 is
   component MultTable_comb_uid191 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid191
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_comb_uid193
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_comb_uid193 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_comb_uid193 is
   component MultTable_comb_uid195 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_comb_uid195
      port map ( X => Xtable,
                 Y => Y1);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_25_comb_uid315
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_25_comb_uid315 is
    port (X : in  std_logic_vector(24 downto 0);
          Y : in  std_logic_vector(24 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(24 downto 0)   );
end entity;

architecture arch of IntAdder_25_comb_uid315 is
signal Rtmp :  std_logic_vector(24 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--       FixMultAdd_signed_x_5_M10_y_5_M10_a_11_M20_r_11_M20_comb_uid2
-- VHDL generated for Kintex7 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan, 2012-2014, 2024
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y A
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixMultAdd_signed_x_5_M10_y_5_M10_a_11_M20_r_11_M20_comb_uid2 is
    port (X : in  std_logic_vector(15 downto 0);
          Y : in  std_logic_vector(15 downto 0);
          A : in  std_logic_vector(31 downto 0);
          R : out  std_logic_vector(31 downto 0)   );
end entity;

architecture arch of FixMultAdd_signed_x_5_M10_y_5_M10_a_11_M20_r_11_M20_comb_uid2 is
   component IntMultiplierLUT_1_signedx2_signed_comb_uid5 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_signed_comb_uid9 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_signed_comb_uid13 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_signed_comb_uid17 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_signed_comb_uid21 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_signed_comb_uid25 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid29 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid33 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid37 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid41 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid45 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid49 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid53 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid57 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid61 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid65 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid69 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid73 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid77 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid81 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid85 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid89 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid93 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid97 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid101 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid105 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid109 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid113 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid117 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid121 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid125 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid129 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid133 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid137 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid141 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid145 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid149 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid153 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid157 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid161 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid165 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid169 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1_signedx2_comb_uid173 is
      port ( X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid177 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid181 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid185 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid189 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_comb_uid193 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_comb_uid198 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_comb_uid201 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_comb_uid204 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_comb_uid209 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_25_comb_uid315 is
      port ( X : in  std_logic_vector(24 downto 0);
             Y : in  std_logic_vector(24 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(24 downto 0)   );
   end component;

signal XX :  signed(5+10 downto 0);
signal YY :  signed(5+10 downto 0);
signal AA :  signed(11+20 downto 0);
signal tile_0_X :  std_logic_vector(0 downto 0);
signal tile_0_Y :  std_logic_vector(1 downto 0);
signal tile_0_output :  std_logic_vector(2 downto 0);
signal tile_0_filtered_output :  signed(2-0 downto 0);
signal bh3_w9_0 :  std_logic;
signal bh3_w10_0 :  std_logic;
signal bh3_w11_0 :  std_logic;
signal tile_1_X :  std_logic_vector(2 downto 0);
signal tile_1_Y :  std_logic_vector(1 downto 0);
signal tile_1_output :  std_logic_vector(4 downto 0);
signal tile_1_filtered_output :  signed(4-0 downto 0);
signal bh3_w6_0 :  std_logic;
signal bh3_w7_0 :  std_logic;
signal bh3_w8_0 :  std_logic;
signal bh3_w9_1 :  std_logic;
signal bh3_w10_1 :  std_logic;
signal tile_2_X :  std_logic_vector(2 downto 0);
signal tile_2_Y :  std_logic_vector(1 downto 0);
signal tile_2_output :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output :  signed(4-0 downto 0);
signal bh3_w3_0 :  std_logic;
signal bh3_w4_0 :  std_logic;
signal bh3_w5_0 :  std_logic;
signal bh3_w6_1 :  std_logic;
signal bh3_w7_1 :  std_logic;
signal tile_3_X :  std_logic_vector(2 downto 0);
signal tile_3_Y :  std_logic_vector(1 downto 0);
signal tile_3_output :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output :  signed(4-0 downto 0);
signal bh3_w0_0 :  std_logic;
signal bh3_w1_0 :  std_logic;
signal bh3_w2_0 :  std_logic;
signal bh3_w3_1 :  std_logic;
signal bh3_w4_1 :  std_logic;
signal tile_4_X :  std_logic_vector(2 downto 0);
signal tile_4_Y :  std_logic_vector(1 downto 0);
signal tile_4_output :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output :  signed(4-0 downto 0);
signal bh3_wm3_0 :  std_logic;
signal bh3_wm2_0 :  std_logic;
signal bh3_wm1_0 :  std_logic;
signal bh3_w0_1 :  std_logic;
signal bh3_w1_1 :  std_logic;
signal tile_5_X :  std_logic_vector(2 downto 0);
signal tile_5_Y :  std_logic_vector(1 downto 0);
signal tile_5_output :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output :  signed(4-0 downto 0);
signal bh3_wm6_0 :  std_logic;
signal bh3_wm5_0 :  std_logic;
signal bh3_wm4_0 :  std_logic;
signal bh3_wm3_1 :  std_logic;
signal bh3_wm2_1 :  std_logic;
signal tile_6_X :  std_logic_vector(0 downto 0);
signal tile_6_Y :  std_logic_vector(1 downto 0);
signal tile_6_output :  std_logic_vector(2 downto 0);
signal tile_6_filtered_output :  signed(2-0 downto 0);
signal bh3_w7_2 :  std_logic;
signal bh3_w8_1 :  std_logic;
signal bh3_w9_2 :  std_logic;
signal tile_7_X :  std_logic_vector(2 downto 0);
signal tile_7_Y :  std_logic_vector(1 downto 0);
signal tile_7_output :  std_logic_vector(4 downto 0);
signal tile_7_filtered_output :  unsigned(4-0 downto 0);
signal bh3_w4_2 :  std_logic;
signal bh3_w5_1 :  std_logic;
signal bh3_w6_2 :  std_logic;
signal bh3_w7_3 :  std_logic;
signal bh3_w8_2 :  std_logic;
signal tile_8_X :  std_logic_vector(2 downto 0);
signal tile_8_Y :  std_logic_vector(1 downto 0);
signal tile_8_output :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output :  unsigned(4-0 downto 0);
signal bh3_w1_2 :  std_logic;
signal bh3_w2_1 :  std_logic;
signal bh3_w3_2 :  std_logic;
signal bh3_w4_3 :  std_logic;
signal bh3_w5_2 :  std_logic;
signal tile_9_X :  std_logic_vector(2 downto 0);
signal tile_9_Y :  std_logic_vector(1 downto 0);
signal tile_9_output :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm2_2 :  std_logic;
signal bh3_wm1_1 :  std_logic;
signal bh3_w0_2 :  std_logic;
signal bh3_w1_3 :  std_logic;
signal bh3_w2_2 :  std_logic;
signal tile_10_X :  std_logic_vector(2 downto 0);
signal tile_10_Y :  std_logic_vector(1 downto 0);
signal tile_10_output :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm5_1 :  std_logic;
signal bh3_wm4_1 :  std_logic;
signal bh3_wm3_2 :  std_logic;
signal bh3_wm2_3 :  std_logic;
signal bh3_wm1_2 :  std_logic;
signal tile_11_X :  std_logic_vector(2 downto 0);
signal tile_11_Y :  std_logic_vector(1 downto 0);
signal tile_11_output :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm8_0 :  std_logic;
signal bh3_wm7_0 :  std_logic;
signal bh3_wm6_1 :  std_logic;
signal bh3_wm5_2 :  std_logic;
signal bh3_wm4_2 :  std_logic;
signal tile_12_X :  std_logic_vector(0 downto 0);
signal tile_12_Y :  std_logic_vector(1 downto 0);
signal tile_12_output :  std_logic_vector(2 downto 0);
signal tile_12_filtered_output :  signed(2-0 downto 0);
signal bh3_w5_3 :  std_logic;
signal bh3_w6_3 :  std_logic;
signal bh3_w7_4 :  std_logic;
signal tile_13_X :  std_logic_vector(2 downto 0);
signal tile_13_Y :  std_logic_vector(1 downto 0);
signal tile_13_output :  std_logic_vector(4 downto 0);
signal tile_13_filtered_output :  unsigned(4-0 downto 0);
signal bh3_w2_3 :  std_logic;
signal bh3_w3_3 :  std_logic;
signal bh3_w4_4 :  std_logic;
signal bh3_w5_4 :  std_logic;
signal bh3_w6_4 :  std_logic;
signal tile_14_X :  std_logic_vector(2 downto 0);
signal tile_14_Y :  std_logic_vector(1 downto 0);
signal tile_14_output :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm1_3 :  std_logic;
signal bh3_w0_3 :  std_logic;
signal bh3_w1_4 :  std_logic;
signal bh3_w2_4 :  std_logic;
signal bh3_w3_4 :  std_logic;
signal tile_15_X :  std_logic_vector(2 downto 0);
signal tile_15_Y :  std_logic_vector(1 downto 0);
signal tile_15_output :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm4_3 :  std_logic;
signal bh3_wm3_3 :  std_logic;
signal bh3_wm2_4 :  std_logic;
signal bh3_wm1_4 :  std_logic;
signal bh3_w0_4 :  std_logic;
signal tile_16_X :  std_logic_vector(2 downto 0);
signal tile_16_Y :  std_logic_vector(1 downto 0);
signal tile_16_output :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm7_1 :  std_logic;
signal bh3_wm6_2 :  std_logic;
signal bh3_wm5_3 :  std_logic;
signal bh3_wm4_4 :  std_logic;
signal bh3_wm3_4 :  std_logic;
signal tile_17_X :  std_logic_vector(2 downto 0);
signal tile_17_Y :  std_logic_vector(1 downto 0);
signal tile_17_output :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm10_0 :  std_logic;
signal bh3_wm9_0 :  std_logic;
signal bh3_wm8_1 :  std_logic;
signal bh3_wm7_2 :  std_logic;
signal bh3_wm6_3 :  std_logic;
signal tile_18_X :  std_logic_vector(0 downto 0);
signal tile_18_Y :  std_logic_vector(1 downto 0);
signal tile_18_output :  std_logic_vector(2 downto 0);
signal tile_18_filtered_output :  signed(2-0 downto 0);
signal bh3_w3_5 :  std_logic;
signal bh3_w4_5 :  std_logic;
signal bh3_w5_5 :  std_logic;
signal tile_19_X :  std_logic_vector(2 downto 0);
signal tile_19_Y :  std_logic_vector(1 downto 0);
signal tile_19_output :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output :  unsigned(4-0 downto 0);
signal bh3_w0_5 :  std_logic;
signal bh3_w1_5 :  std_logic;
signal bh3_w2_5 :  std_logic;
signal bh3_w3_6 :  std_logic;
signal bh3_w4_6 :  std_logic;
signal tile_20_X :  std_logic_vector(2 downto 0);
signal tile_20_Y :  std_logic_vector(1 downto 0);
signal tile_20_output :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm3_5 :  std_logic;
signal bh3_wm2_5 :  std_logic;
signal bh3_wm1_5 :  std_logic;
signal bh3_w0_6 :  std_logic;
signal bh3_w1_6 :  std_logic;
signal tile_21_X :  std_logic_vector(2 downto 0);
signal tile_21_Y :  std_logic_vector(1 downto 0);
signal tile_21_output :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm6_4 :  std_logic;
signal bh3_wm5_4 :  std_logic;
signal bh3_wm4_5 :  std_logic;
signal bh3_wm3_6 :  std_logic;
signal bh3_wm2_6 :  std_logic;
signal tile_22_X :  std_logic_vector(2 downto 0);
signal tile_22_Y :  std_logic_vector(1 downto 0);
signal tile_22_output :  std_logic_vector(4 downto 0);
signal tile_22_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm9_1 :  std_logic;
signal bh3_wm8_2 :  std_logic;
signal bh3_wm7_3 :  std_logic;
signal bh3_wm6_5 :  std_logic;
signal bh3_wm5_5 :  std_logic;
signal tile_23_X :  std_logic_vector(2 downto 0);
signal tile_23_Y :  std_logic_vector(1 downto 0);
signal tile_23_output :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm12_0 :  std_logic;
signal bh3_wm11_0 :  std_logic;
signal bh3_wm10_1 :  std_logic;
signal bh3_wm9_2 :  std_logic;
signal bh3_wm8_3 :  std_logic;
signal tile_24_X :  std_logic_vector(0 downto 0);
signal tile_24_Y :  std_logic_vector(1 downto 0);
signal tile_24_output :  std_logic_vector(2 downto 0);
signal tile_24_filtered_output :  signed(2-0 downto 0);
signal bh3_w1_7 :  std_logic;
signal bh3_w2_6 :  std_logic;
signal bh3_w3_7 :  std_logic;
signal tile_25_X :  std_logic_vector(2 downto 0);
signal tile_25_Y :  std_logic_vector(1 downto 0);
signal tile_25_output :  std_logic_vector(4 downto 0);
signal tile_25_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm2_7 :  std_logic;
signal bh3_wm1_6 :  std_logic;
signal bh3_w0_7 :  std_logic;
signal bh3_w1_8 :  std_logic;
signal bh3_w2_7 :  std_logic;
signal tile_26_X :  std_logic_vector(2 downto 0);
signal tile_26_Y :  std_logic_vector(1 downto 0);
signal tile_26_output :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm5_6 :  std_logic;
signal bh3_wm4_6 :  std_logic;
signal bh3_wm3_7 :  std_logic;
signal bh3_wm2_8 :  std_logic;
signal bh3_wm1_7 :  std_logic;
signal tile_27_X :  std_logic_vector(2 downto 0);
signal tile_27_Y :  std_logic_vector(1 downto 0);
signal tile_27_output :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm8_4 :  std_logic;
signal bh3_wm7_4 :  std_logic;
signal bh3_wm6_6 :  std_logic;
signal bh3_wm5_7 :  std_logic;
signal bh3_wm4_7 :  std_logic;
signal tile_28_X :  std_logic_vector(2 downto 0);
signal tile_28_Y :  std_logic_vector(1 downto 0);
signal tile_28_output :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm11_1 :  std_logic;
signal bh3_wm10_2 :  std_logic;
signal bh3_wm9_3 :  std_logic;
signal bh3_wm8_5 :  std_logic;
signal bh3_wm7_5 :  std_logic;
signal tile_29_X :  std_logic_vector(2 downto 0);
signal tile_29_Y :  std_logic_vector(1 downto 0);
signal tile_29_output :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm14_0 :  std_logic;
signal bh3_wm13_0 :  std_logic;
signal bh3_wm12_1 :  std_logic;
signal bh3_wm11_2 :  std_logic;
signal bh3_wm10_3 :  std_logic;
signal tile_30_X :  std_logic_vector(0 downto 0);
signal tile_30_Y :  std_logic_vector(1 downto 0);
signal tile_30_output :  std_logic_vector(2 downto 0);
signal tile_30_filtered_output :  signed(2-0 downto 0);
signal bh3_wm1_8 :  std_logic;
signal bh3_w0_8 :  std_logic;
signal bh3_w1_9 :  std_logic;
signal tile_31_X :  std_logic_vector(2 downto 0);
signal tile_31_Y :  std_logic_vector(1 downto 0);
signal tile_31_output :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm4_8 :  std_logic;
signal bh3_wm3_8 :  std_logic;
signal bh3_wm2_9 :  std_logic;
signal bh3_wm1_9 :  std_logic;
signal bh3_w0_9 :  std_logic;
signal tile_32_X :  std_logic_vector(2 downto 0);
signal tile_32_Y :  std_logic_vector(1 downto 0);
signal tile_32_output :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm7_6 :  std_logic;
signal bh3_wm6_7 :  std_logic;
signal bh3_wm5_8 :  std_logic;
signal bh3_wm4_9 :  std_logic;
signal bh3_wm3_9 :  std_logic;
signal tile_33_X :  std_logic_vector(2 downto 0);
signal tile_33_Y :  std_logic_vector(1 downto 0);
signal tile_33_output :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm10_4 :  std_logic;
signal bh3_wm9_4 :  std_logic;
signal bh3_wm8_6 :  std_logic;
signal bh3_wm7_7 :  std_logic;
signal bh3_wm6_8 :  std_logic;
signal tile_34_X :  std_logic_vector(2 downto 0);
signal tile_34_Y :  std_logic_vector(1 downto 0);
signal tile_34_output :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm13_1 :  std_logic;
signal bh3_wm12_2 :  std_logic;
signal bh3_wm11_3 :  std_logic;
signal bh3_wm10_5 :  std_logic;
signal bh3_wm9_5 :  std_logic;
signal tile_35_X :  std_logic_vector(2 downto 0);
signal tile_35_Y :  std_logic_vector(1 downto 0);
signal tile_35_output :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm16_0 :  std_logic;
signal bh3_wm15_0 :  std_logic;
signal bh3_wm14_1 :  std_logic;
signal bh3_wm13_2 :  std_logic;
signal bh3_wm12_3 :  std_logic;
signal tile_36_X :  std_logic_vector(0 downto 0);
signal tile_36_Y :  std_logic_vector(1 downto 0);
signal tile_36_output :  std_logic_vector(2 downto 0);
signal tile_36_filtered_output :  signed(2-0 downto 0);
signal bh3_wm3_10 :  std_logic;
signal bh3_wm2_10 :  std_logic;
signal bh3_wm1_10 :  std_logic;
signal tile_37_X :  std_logic_vector(2 downto 0);
signal tile_37_Y :  std_logic_vector(1 downto 0);
signal tile_37_output :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm6_9 :  std_logic;
signal bh3_wm5_9 :  std_logic;
signal bh3_wm4_10 :  std_logic;
signal bh3_wm3_11 :  std_logic;
signal bh3_wm2_11 :  std_logic;
signal tile_38_X :  std_logic_vector(2 downto 0);
signal tile_38_Y :  std_logic_vector(1 downto 0);
signal tile_38_output :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm9_6 :  std_logic;
signal bh3_wm8_7 :  std_logic;
signal bh3_wm7_8 :  std_logic;
signal bh3_wm6_10 :  std_logic;
signal bh3_wm5_10 :  std_logic;
signal tile_39_X :  std_logic_vector(2 downto 0);
signal tile_39_Y :  std_logic_vector(1 downto 0);
signal tile_39_output :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm12_4 :  std_logic;
signal bh3_wm11_4 :  std_logic;
signal bh3_wm10_6 :  std_logic;
signal bh3_wm9_7 :  std_logic;
signal bh3_wm8_8 :  std_logic;
signal tile_40_X :  std_logic_vector(2 downto 0);
signal tile_40_Y :  std_logic_vector(1 downto 0);
signal tile_40_output :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm15_1 :  std_logic;
signal bh3_wm14_2 :  std_logic;
signal bh3_wm13_3 :  std_logic;
signal bh3_wm12_5 :  std_logic;
signal bh3_wm11_5 :  std_logic;
signal tile_41_X :  std_logic_vector(2 downto 0);
signal tile_41_Y :  std_logic_vector(1 downto 0);
signal tile_41_output :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm18_0 :  std_logic;
signal bh3_wm17_0 :  std_logic;
signal bh3_wm16_1 :  std_logic;
signal bh3_wm15_2 :  std_logic;
signal bh3_wm14_3 :  std_logic;
signal tile_42_X :  std_logic_vector(0 downto 0);
signal tile_42_Y :  std_logic_vector(1 downto 0);
signal tile_42_output :  std_logic_vector(2 downto 0);
signal tile_42_filtered_output :  signed(2-0 downto 0);
signal bh3_wm5_11 :  std_logic;
signal bh3_wm4_11 :  std_logic;
signal bh3_wm3_12 :  std_logic;
signal tile_43_X :  std_logic_vector(2 downto 0);
signal tile_43_Y :  std_logic_vector(1 downto 0);
signal tile_43_output :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm8_9 :  std_logic;
signal bh3_wm7_9 :  std_logic;
signal bh3_wm6_11 :  std_logic;
signal bh3_wm5_12 :  std_logic;
signal bh3_wm4_12 :  std_logic;
signal tile_44_X :  std_logic_vector(2 downto 0);
signal tile_44_Y :  std_logic_vector(1 downto 0);
signal tile_44_output :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm11_6 :  std_logic;
signal bh3_wm10_7 :  std_logic;
signal bh3_wm9_8 :  std_logic;
signal bh3_wm8_10 :  std_logic;
signal bh3_wm7_10 :  std_logic;
signal tile_45_X :  std_logic_vector(2 downto 0);
signal tile_45_Y :  std_logic_vector(1 downto 0);
signal tile_45_output :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm14_4 :  std_logic;
signal bh3_wm13_4 :  std_logic;
signal bh3_wm12_6 :  std_logic;
signal bh3_wm11_7 :  std_logic;
signal bh3_wm10_8 :  std_logic;
signal tile_46_X :  std_logic_vector(2 downto 0);
signal tile_46_Y :  std_logic_vector(1 downto 0);
signal tile_46_output :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm17_1 :  std_logic;
signal bh3_wm16_2 :  std_logic;
signal bh3_wm15_3 :  std_logic;
signal bh3_wm14_5 :  std_logic;
signal bh3_wm13_5 :  std_logic;
signal tile_47_X :  std_logic_vector(2 downto 0);
signal tile_47_Y :  std_logic_vector(1 downto 0);
signal tile_47_output :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output :  unsigned(4-0 downto 0);
signal bh3_wm20_0 :  std_logic;
signal bh3_wm19_0 :  std_logic;
signal bh3_wm18_1 :  std_logic;
signal bh3_wm17_2 :  std_logic;
signal bh3_wm16_3 :  std_logic;
signal bh3_wm20_1 :  std_logic;
signal bh3_wm19_1 :  std_logic;
signal bh3_wm18_2 :  std_logic;
signal bh3_wm17_3 :  std_logic;
signal bh3_wm16_4 :  std_logic;
signal bh3_wm15_4 :  std_logic;
signal bh3_wm14_6 :  std_logic;
signal bh3_wm13_6 :  std_logic;
signal bh3_wm12_7 :  std_logic;
signal bh3_wm11_8 :  std_logic;
signal bh3_wm10_9 :  std_logic;
signal bh3_wm9_9 :  std_logic;
signal bh3_wm8_11 :  std_logic;
signal bh3_wm7_11 :  std_logic;
signal bh3_wm6_12 :  std_logic;
signal bh3_wm5_13 :  std_logic;
signal bh3_wm4_13 :  std_logic;
signal bh3_wm3_13 :  std_logic;
signal bh3_wm2_12 :  std_logic;
signal bh3_wm1_11 :  std_logic;
signal bh3_w0_10 :  std_logic;
signal bh3_w1_10 :  std_logic;
signal bh3_w2_8 :  std_logic;
signal bh3_w3_8 :  std_logic;
signal bh3_w4_7 :  std_logic;
signal bh3_w5_6 :  std_logic;
signal bh3_w6_5 :  std_logic;
signal bh3_w7_5 :  std_logic;
signal bh3_w8_3 :  std_logic;
signal bh3_w9_3 :  std_logic;
signal bh3_w10_2 :  std_logic;
signal bh3_w11_1 :  std_logic;
signal bh3_wm3_14 :  std_logic;
signal bh3_w0_11 :  std_logic;
signal bh3_w1_11 :  std_logic;
signal bh3_w6_6 :  std_logic;
signal bh3_w7_6 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid199_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid199_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid199_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm20_2 :  std_logic;
signal bh3_wm19_2 :  std_logic;
signal bh3_wm18_3 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid202_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid202_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm18_4 :  std_logic;
signal bh3_wm17_4 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid205_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid205_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid205_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm17_5 :  std_logic;
signal bh3_wm16_5 :  std_logic;
signal bh3_wm15_5 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid206_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid206_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid206_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm16_6 :  std_logic;
signal bh3_wm15_6 :  std_logic;
signal bh3_wm14_7 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid207_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid207_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid207_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm15_7 :  std_logic;
signal bh3_wm14_8 :  std_logic;
signal bh3_wm13_7 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid210_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid210_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm14_9 :  std_logic;
signal bh3_wm13_8 :  std_logic;
signal bh3_wm12_8 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid211_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid211_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm13_9 :  std_logic;
signal bh3_wm12_9 :  std_logic;
signal bh3_wm11_9 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid212_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid212_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid212_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm13_10 :  std_logic;
signal bh3_wm12_10 :  std_logic;
signal bh3_wm11_10 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid213_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid213_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm12_11 :  std_logic;
signal bh3_wm11_11 :  std_logic;
signal bh3_wm10_10 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid214_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid214_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm11_12 :  std_logic;
signal bh3_wm10_11 :  std_logic;
signal bh3_wm9_10 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid215_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid215_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm11_13 :  std_logic;
signal bh3_wm10_12 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid216_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid216_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm10_13 :  std_logic;
signal bh3_wm9_11 :  std_logic;
signal bh3_wm8_12 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid217_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid217_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid217_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm10_14 :  std_logic;
signal bh3_wm9_12 :  std_logic;
signal bh3_wm8_13 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid218_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid218_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm9_13 :  std_logic;
signal bh3_wm8_14 :  std_logic;
signal bh3_wm7_12 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid219_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid219_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm9_14 :  std_logic;
signal bh3_wm8_15 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid220_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid220_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm8_16 :  std_logic;
signal bh3_wm7_13 :  std_logic;
signal bh3_wm6_13 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid221_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid221_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm8_17 :  std_logic;
signal bh3_wm7_14 :  std_logic;
signal bh3_wm6_14 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid222_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid222_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm7_15 :  std_logic;
signal bh3_wm6_15 :  std_logic;
signal bh3_wm5_14 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid223_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid223_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm7_16 :  std_logic;
signal bh3_wm6_16 :  std_logic;
signal bh3_wm5_15 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid224_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid224_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm6_17 :  std_logic;
signal bh3_wm5_16 :  std_logic;
signal bh3_wm4_14 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid225_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid225_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm6_18 :  std_logic;
signal bh3_wm5_17 :  std_logic;
signal bh3_wm4_15 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid226_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid226_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm5_18 :  std_logic;
signal bh3_wm4_16 :  std_logic;
signal bh3_wm3_15 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid227_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid227_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm5_19 :  std_logic;
signal bh3_wm4_17 :  std_logic;
signal bh3_wm3_16 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid228_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid228_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid228_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm5_20 :  std_logic;
signal bh3_wm4_18 :  std_logic;
signal bh3_wm3_17 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid229_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid229_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm4_19 :  std_logic;
signal bh3_wm3_18 :  std_logic;
signal bh3_wm2_13 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid230_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid230_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm4_20 :  std_logic;
signal bh3_wm3_19 :  std_logic;
signal bh3_wm2_14 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid231_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid231_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm3_20 :  std_logic;
signal bh3_wm2_15 :  std_logic;
signal bh3_wm1_12 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid232_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid232_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm3_21 :  std_logic;
signal bh3_wm2_16 :  std_logic;
signal bh3_wm1_13 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid233_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid233_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm3_22 :  std_logic;
signal bh3_wm2_17 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid234_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid234_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm2_18 :  std_logic;
signal bh3_wm1_14 :  std_logic;
signal bh3_w0_12 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid235_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid235_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm2_19 :  std_logic;
signal bh3_wm1_15 :  std_logic;
signal bh3_w0_13 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid236_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid236_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm1_16 :  std_logic;
signal bh3_w0_14 :  std_logic;
signal bh3_w1_12 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid237_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid237_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm1_17 :  std_logic;
signal bh3_w0_15 :  std_logic;
signal bh3_w1_13 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid238_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid238_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w0_16 :  std_logic;
signal bh3_w1_14 :  std_logic;
signal bh3_w2_9 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid239_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid239_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w0_17 :  std_logic;
signal bh3_w1_15 :  std_logic;
signal bh3_w2_10 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid240_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid240_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w1_16 :  std_logic;
signal bh3_w2_11 :  std_logic;
signal bh3_w3_9 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid241_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid241_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w1_17 :  std_logic;
signal bh3_w2_12 :  std_logic;
signal bh3_w3_10 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid242_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid242_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w2_13 :  std_logic;
signal bh3_w3_11 :  std_logic;
signal bh3_w4_8 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid243_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid243_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid243_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w2_14 :  std_logic;
signal bh3_w3_12 :  std_logic;
signal bh3_w4_9 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid244_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid244_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w3_13 :  std_logic;
signal bh3_w4_10 :  std_logic;
signal bh3_w5_7 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid245_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid245_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w4_11 :  std_logic;
signal bh3_w5_8 :  std_logic;
signal bh3_w6_7 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid246_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid246_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid246_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w4_12 :  std_logic;
signal bh3_w5_9 :  std_logic;
signal bh3_w6_8 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid247_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid247_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w5_10 :  std_logic;
signal bh3_w6_9 :  std_logic;
signal bh3_w7_7 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid248_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid248_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w6_10 :  std_logic;
signal bh3_w7_8 :  std_logic;
signal bh3_w8_4 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid249_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid249_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w7_9 :  std_logic;
signal bh3_w8_5 :  std_logic;
signal bh3_w9_4 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid250_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid250_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid250_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w8_6 :  std_logic;
signal bh3_w9_5 :  std_logic;
signal bh3_w10_3 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid251_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid251_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid251_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w9_6 :  std_logic;
signal bh3_w10_4 :  std_logic;
signal bh3_w11_2 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid252_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid252_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid252_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w10_5 :  std_logic;
signal bh3_w11_3 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid253_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid253_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid253_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm18_5 :  std_logic;
signal bh3_wm17_6 :  std_logic;
signal bh3_wm16_7 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid254_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid254_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm16_8 :  std_logic;
signal bh3_wm15_8 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid255_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid255_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid255_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm15_9 :  std_logic;
signal bh3_wm14_10 :  std_logic;
signal bh3_wm13_11 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid256_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid256_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid256_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm13_12 :  std_logic;
signal bh3_wm12_12 :  std_logic;
signal bh3_wm11_14 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid257_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid257_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm12_13 :  std_logic;
signal bh3_wm11_15 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid258_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid258_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid258_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm11_16 :  std_logic;
signal bh3_wm10_15 :  std_logic;
signal bh3_wm9_15 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid259_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid259_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid259_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm10_16 :  std_logic;
signal bh3_wm9_16 :  std_logic;
signal bh3_wm8_18 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid260_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid260_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm9_17 :  std_logic;
signal bh3_wm8_19 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid261_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid261_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm8_20 :  std_logic;
signal bh3_wm7_17 :  std_logic;
signal bh3_wm6_19 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid262_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid262_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid262_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm7_18 :  std_logic;
signal bh3_wm6_20 :  std_logic;
signal bh3_wm5_21 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid263_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid263_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm6_21 :  std_logic;
signal bh3_wm5_22 :  std_logic;
signal bh3_wm4_21 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid264_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid264_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm5_23 :  std_logic;
signal bh3_wm4_22 :  std_logic;
signal bh3_wm3_23 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid265_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid265_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm4_23 :  std_logic;
signal bh3_wm3_24 :  std_logic;
signal bh3_wm2_20 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid266_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid266_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm3_25 :  std_logic;
signal bh3_wm2_21 :  std_logic;
signal bh3_wm1_18 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid267_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid267_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid267_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm3_26 :  std_logic;
signal bh3_wm2_22 :  std_logic;
signal bh3_wm1_19 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid268_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid268_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm2_23 :  std_logic;
signal bh3_wm1_20 :  std_logic;
signal bh3_w0_18 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid269_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid269_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm1_21 :  std_logic;
signal bh3_w0_19 :  std_logic;
signal bh3_w1_18 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid270_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid270_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w0_20 :  std_logic;
signal bh3_w1_19 :  std_logic;
signal bh3_w2_15 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid271_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid271_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w1_20 :  std_logic;
signal bh3_w2_16 :  std_logic;
signal bh3_w3_14 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid272_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid272_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w2_17 :  std_logic;
signal bh3_w3_15 :  std_logic;
signal bh3_w4_13 :  std_logic;
signal Compressor_6_3_comb_uid209_bh3_uid273_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_comb_uid209_bh3_uid273_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w3_16 :  std_logic;
signal bh3_w4_14 :  std_logic;
signal bh3_w5_11 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid274_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid274_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid274_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w4_15 :  std_logic;
signal bh3_w5_12 :  std_logic;
signal bh3_w6_11 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid275_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid275_Out0 :  std_logic_vector(1 downto 0);
signal bh3_w5_13 :  std_logic;
signal bh3_w6_12 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid276_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid276_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid276_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w6_13 :  std_logic;
signal bh3_w7_10 :  std_logic;
signal bh3_w8_7 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid277_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid277_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid277_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w7_11 :  std_logic;
signal bh3_w8_8 :  std_logic;
signal bh3_w9_7 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid278_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid278_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid278_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w9_8 :  std_logic;
signal bh3_w10_6 :  std_logic;
signal bh3_w11_4 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid279_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid279_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid279_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w11_5 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid280_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid280_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid280_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm16_9 :  std_logic;
signal bh3_wm15_10 :  std_logic;
signal bh3_wm14_11 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid281_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid281_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid281_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm14_12 :  std_logic;
signal bh3_wm13_13 :  std_logic;
signal bh3_wm12_14 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid282_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid282_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm12_15 :  std_logic;
signal bh3_wm11_17 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid283_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid283_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid283_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm11_18 :  std_logic;
signal bh3_wm10_17 :  std_logic;
signal bh3_wm9_18 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid284_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid284_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid284_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm9_19 :  std_logic;
signal bh3_wm8_21 :  std_logic;
signal bh3_wm7_19 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid285_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid285_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm8_22 :  std_logic;
signal bh3_wm7_20 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid286_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid286_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid286_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm7_21 :  std_logic;
signal bh3_wm6_22 :  std_logic;
signal bh3_wm5_24 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid287_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid287_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid287_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm5_25 :  std_logic;
signal bh3_wm4_24 :  std_logic;
signal bh3_wm3_27 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid288_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid288_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm4_25 :  std_logic;
signal bh3_wm3_28 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid289_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid289_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid289_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm3_29 :  std_logic;
signal bh3_wm2_24 :  std_logic;
signal bh3_wm1_22 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid290_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid290_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm2_25 :  std_logic;
signal bh3_wm1_23 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid291_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid291_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid291_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm1_24 :  std_logic;
signal bh3_w0_21 :  std_logic;
signal bh3_w1_21 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid292_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid292_Out0 :  std_logic_vector(1 downto 0);
signal bh3_w0_22 :  std_logic;
signal bh3_w1_22 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid293_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid293_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid293_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w1_23 :  std_logic;
signal bh3_w2_18 :  std_logic;
signal bh3_w3_17 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid294_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid294_Out0 :  std_logic_vector(1 downto 0);
signal bh3_w3_18 :  std_logic;
signal bh3_w4_16 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid295_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid295_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid295_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w4_17 :  std_logic;
signal bh3_w5_14 :  std_logic;
signal bh3_w6_14 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid296_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid296_Out0 :  std_logic_vector(1 downto 0);
signal bh3_w5_15 :  std_logic;
signal bh3_w6_15 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid297_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid297_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid297_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w6_16 :  std_logic;
signal bh3_w7_12 :  std_logic;
signal bh3_w8_9 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid298_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid298_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid298_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w8_10 :  std_logic;
signal bh3_w9_9 :  std_logic;
signal bh3_w10_7 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid299_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid299_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid299_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w10_8 :  std_logic;
signal bh3_w11_6 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid300_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid300_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid300_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm14_13 :  std_logic;
signal bh3_wm13_14 :  std_logic;
signal bh3_wm12_16 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid301_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid301_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid301_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm12_17 :  std_logic;
signal bh3_wm11_19 :  std_logic;
signal bh3_wm10_18 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid302_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid302_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid302_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm10_19 :  std_logic;
signal bh3_wm9_20 :  std_logic;
signal bh3_wm8_23 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid303_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid303_Out0 :  std_logic_vector(1 downto 0);
signal bh3_wm8_24 :  std_logic;
signal bh3_wm7_22 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid304_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid304_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid304_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm7_23 :  std_logic;
signal bh3_wm6_23 :  std_logic;
signal bh3_wm5_26 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid305_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid305_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid305_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm5_27 :  std_logic;
signal bh3_wm4_26 :  std_logic;
signal bh3_wm3_30 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid306_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid306_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid306_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm3_31 :  std_logic;
signal bh3_wm2_26 :  std_logic;
signal bh3_wm1_25 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid307_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid307_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid307_Out0 :  std_logic_vector(2 downto 0);
signal bh3_wm1_26 :  std_logic;
signal bh3_w0_23 :  std_logic;
signal bh3_w1_24 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid308_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid308_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid308_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w1_25 :  std_logic;
signal bh3_w2_19 :  std_logic;
signal bh3_w3_19 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid309_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid309_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid309_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w3_20 :  std_logic;
signal bh3_w4_18 :  std_logic;
signal bh3_w5_16 :  std_logic;
signal Compressor_3_2_comb_uid201_bh3_uid310_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_comb_uid201_bh3_uid310_Out0 :  std_logic_vector(1 downto 0);
signal bh3_w5_17 :  std_logic;
signal bh3_w6_17 :  std_logic;
signal Compressor_23_3_comb_uid198_bh3_uid311_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid311_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_comb_uid198_bh3_uid311_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w6_18 :  std_logic;
signal bh3_w7_13 :  std_logic;
signal bh3_w8_11 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid312_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid312_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid312_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w8_12 :  std_logic;
signal bh3_w9_10 :  std_logic;
signal bh3_w10_9 :  std_logic;
signal Compressor_14_3_comb_uid204_bh3_uid313_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid313_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_comb_uid204_bh3_uid313_Out0 :  std_logic_vector(2 downto 0);
signal bh3_w10_10 :  std_logic;
signal bh3_w11_7 :  std_logic;
signal tmp_bitheapResult_bh3_7 :  std_logic_vector(7 downto 0);
signal bitheapFinalAdd_bh3_In0 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh3_In1 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh3_Cin :  std_logic;
signal bitheapFinalAdd_bh3_Out :  std_logic_vector(24 downto 0);
signal bitheapResult_bh3 :  std_logic_vector(31 downto 0);
signal RR :  signed(11+20 downto 0);
begin
XX <= signed(X);
YY <= signed(Y);
AA <= signed(A);
   tile_0_X <= X(15 downto 15);
   tile_0_Y <= Y(15 downto 14);
   tile_0_mult: IntMultiplierLUT_1_signedx2_signed_comb_uid5
      port map ( X => tile_0_X,
                 Y => tile_0_Y,
                 R => tile_0_output);

   tile_0_filtered_output <= signed(tile_0_output(2 downto 0));
   bh3_w9_0 <= tile_0_filtered_output(0);
   bh3_w10_0 <= tile_0_filtered_output(1);
   bh3_w11_0 <= not tile_0_filtered_output(2);
   tile_1_X <= X(14 downto 12);
   tile_1_Y <= Y(15 downto 14);
   tile_1_mult: IntMultiplierLUT_3x2_signed_comb_uid9
      port map ( X => tile_1_X,
                 Y => tile_1_Y,
                 R => tile_1_output);

   tile_1_filtered_output <= signed(tile_1_output(4 downto 0));
   bh3_w6_0 <= tile_1_filtered_output(0);
   bh3_w7_0 <= tile_1_filtered_output(1);
   bh3_w8_0 <= tile_1_filtered_output(2);
   bh3_w9_1 <= tile_1_filtered_output(3);
   bh3_w10_1 <= not tile_1_filtered_output(4);
   tile_2_X <= X(11 downto 9);
   tile_2_Y <= Y(15 downto 14);
   tile_2_mult: IntMultiplierLUT_3x2_signed_comb_uid13
      port map ( X => tile_2_X,
                 Y => tile_2_Y,
                 R => tile_2_output);

   tile_2_filtered_output <= signed(tile_2_output(4 downto 0));
   bh3_w3_0 <= tile_2_filtered_output(0);
   bh3_w4_0 <= tile_2_filtered_output(1);
   bh3_w5_0 <= tile_2_filtered_output(2);
   bh3_w6_1 <= tile_2_filtered_output(3);
   bh3_w7_1 <= not tile_2_filtered_output(4);
   tile_3_X <= X(8 downto 6);
   tile_3_Y <= Y(15 downto 14);
   tile_3_mult: IntMultiplierLUT_3x2_signed_comb_uid17
      port map ( X => tile_3_X,
                 Y => tile_3_Y,
                 R => tile_3_output);

   tile_3_filtered_output <= signed(tile_3_output(4 downto 0));
   bh3_w0_0 <= tile_3_filtered_output(0);
   bh3_w1_0 <= tile_3_filtered_output(1);
   bh3_w2_0 <= tile_3_filtered_output(2);
   bh3_w3_1 <= tile_3_filtered_output(3);
   bh3_w4_1 <= not tile_3_filtered_output(4);
   tile_4_X <= X(5 downto 3);
   tile_4_Y <= Y(15 downto 14);
   tile_4_mult: IntMultiplierLUT_3x2_signed_comb_uid21
      port map ( X => tile_4_X,
                 Y => tile_4_Y,
                 R => tile_4_output);

   tile_4_filtered_output <= signed(tile_4_output(4 downto 0));
   bh3_wm3_0 <= tile_4_filtered_output(0);
   bh3_wm2_0 <= tile_4_filtered_output(1);
   bh3_wm1_0 <= tile_4_filtered_output(2);
   bh3_w0_1 <= tile_4_filtered_output(3);
   bh3_w1_1 <= not tile_4_filtered_output(4);
   tile_5_X <= X(2 downto 0);
   tile_5_Y <= Y(15 downto 14);
   tile_5_mult: IntMultiplierLUT_3x2_signed_comb_uid25
      port map ( X => tile_5_X,
                 Y => tile_5_Y,
                 R => tile_5_output);

   tile_5_filtered_output <= signed(tile_5_output(4 downto 0));
   bh3_wm6_0 <= tile_5_filtered_output(0);
   bh3_wm5_0 <= tile_5_filtered_output(1);
   bh3_wm4_0 <= tile_5_filtered_output(2);
   bh3_wm3_1 <= tile_5_filtered_output(3);
   bh3_wm2_1 <= not tile_5_filtered_output(4);
   tile_6_X <= X(15 downto 15);
   tile_6_Y <= Y(13 downto 12);
   tile_6_mult: IntMultiplierLUT_1_signedx2_comb_uid29
      port map ( X => tile_6_X,
                 Y => tile_6_Y,
                 R => tile_6_output);

   tile_6_filtered_output <= signed(tile_6_output(2 downto 0));
   bh3_w7_2 <= tile_6_filtered_output(0);
   bh3_w8_1 <= tile_6_filtered_output(1);
   bh3_w9_2 <= not tile_6_filtered_output(2);
   tile_7_X <= X(14 downto 12);
   tile_7_Y <= Y(13 downto 12);
   tile_7_mult: IntMultiplierLUT_3x2_comb_uid33
      port map ( X => tile_7_X,
                 Y => tile_7_Y,
                 R => tile_7_output);

   tile_7_filtered_output <= unsigned(tile_7_output(4 downto 0));
   bh3_w4_2 <= tile_7_filtered_output(0);
   bh3_w5_1 <= tile_7_filtered_output(1);
   bh3_w6_2 <= tile_7_filtered_output(2);
   bh3_w7_3 <= tile_7_filtered_output(3);
   bh3_w8_2 <= tile_7_filtered_output(4);
   tile_8_X <= X(11 downto 9);
   tile_8_Y <= Y(13 downto 12);
   tile_8_mult: IntMultiplierLUT_3x2_comb_uid37
      port map ( X => tile_8_X,
                 Y => tile_8_Y,
                 R => tile_8_output);

   tile_8_filtered_output <= unsigned(tile_8_output(4 downto 0));
   bh3_w1_2 <= tile_8_filtered_output(0);
   bh3_w2_1 <= tile_8_filtered_output(1);
   bh3_w3_2 <= tile_8_filtered_output(2);
   bh3_w4_3 <= tile_8_filtered_output(3);
   bh3_w5_2 <= tile_8_filtered_output(4);
   tile_9_X <= X(8 downto 6);
   tile_9_Y <= Y(13 downto 12);
   tile_9_mult: IntMultiplierLUT_3x2_comb_uid41
      port map ( X => tile_9_X,
                 Y => tile_9_Y,
                 R => tile_9_output);

   tile_9_filtered_output <= unsigned(tile_9_output(4 downto 0));
   bh3_wm2_2 <= tile_9_filtered_output(0);
   bh3_wm1_1 <= tile_9_filtered_output(1);
   bh3_w0_2 <= tile_9_filtered_output(2);
   bh3_w1_3 <= tile_9_filtered_output(3);
   bh3_w2_2 <= tile_9_filtered_output(4);
   tile_10_X <= X(5 downto 3);
   tile_10_Y <= Y(13 downto 12);
   tile_10_mult: IntMultiplierLUT_3x2_comb_uid45
      port map ( X => tile_10_X,
                 Y => tile_10_Y,
                 R => tile_10_output);

   tile_10_filtered_output <= unsigned(tile_10_output(4 downto 0));
   bh3_wm5_1 <= tile_10_filtered_output(0);
   bh3_wm4_1 <= tile_10_filtered_output(1);
   bh3_wm3_2 <= tile_10_filtered_output(2);
   bh3_wm2_3 <= tile_10_filtered_output(3);
   bh3_wm1_2 <= tile_10_filtered_output(4);
   tile_11_X <= X(2 downto 0);
   tile_11_Y <= Y(13 downto 12);
   tile_11_mult: IntMultiplierLUT_3x2_comb_uid49
      port map ( X => tile_11_X,
                 Y => tile_11_Y,
                 R => tile_11_output);

   tile_11_filtered_output <= unsigned(tile_11_output(4 downto 0));
   bh3_wm8_0 <= tile_11_filtered_output(0);
   bh3_wm7_0 <= tile_11_filtered_output(1);
   bh3_wm6_1 <= tile_11_filtered_output(2);
   bh3_wm5_2 <= tile_11_filtered_output(3);
   bh3_wm4_2 <= tile_11_filtered_output(4);
   tile_12_X <= X(15 downto 15);
   tile_12_Y <= Y(11 downto 10);
   tile_12_mult: IntMultiplierLUT_1_signedx2_comb_uid53
      port map ( X => tile_12_X,
                 Y => tile_12_Y,
                 R => tile_12_output);

   tile_12_filtered_output <= signed(tile_12_output(2 downto 0));
   bh3_w5_3 <= tile_12_filtered_output(0);
   bh3_w6_3 <= tile_12_filtered_output(1);
   bh3_w7_4 <= not tile_12_filtered_output(2);
   tile_13_X <= X(14 downto 12);
   tile_13_Y <= Y(11 downto 10);
   tile_13_mult: IntMultiplierLUT_3x2_comb_uid57
      port map ( X => tile_13_X,
                 Y => tile_13_Y,
                 R => tile_13_output);

   tile_13_filtered_output <= unsigned(tile_13_output(4 downto 0));
   bh3_w2_3 <= tile_13_filtered_output(0);
   bh3_w3_3 <= tile_13_filtered_output(1);
   bh3_w4_4 <= tile_13_filtered_output(2);
   bh3_w5_4 <= tile_13_filtered_output(3);
   bh3_w6_4 <= tile_13_filtered_output(4);
   tile_14_X <= X(11 downto 9);
   tile_14_Y <= Y(11 downto 10);
   tile_14_mult: IntMultiplierLUT_3x2_comb_uid61
      port map ( X => tile_14_X,
                 Y => tile_14_Y,
                 R => tile_14_output);

   tile_14_filtered_output <= unsigned(tile_14_output(4 downto 0));
   bh3_wm1_3 <= tile_14_filtered_output(0);
   bh3_w0_3 <= tile_14_filtered_output(1);
   bh3_w1_4 <= tile_14_filtered_output(2);
   bh3_w2_4 <= tile_14_filtered_output(3);
   bh3_w3_4 <= tile_14_filtered_output(4);
   tile_15_X <= X(8 downto 6);
   tile_15_Y <= Y(11 downto 10);
   tile_15_mult: IntMultiplierLUT_3x2_comb_uid65
      port map ( X => tile_15_X,
                 Y => tile_15_Y,
                 R => tile_15_output);

   tile_15_filtered_output <= unsigned(tile_15_output(4 downto 0));
   bh3_wm4_3 <= tile_15_filtered_output(0);
   bh3_wm3_3 <= tile_15_filtered_output(1);
   bh3_wm2_4 <= tile_15_filtered_output(2);
   bh3_wm1_4 <= tile_15_filtered_output(3);
   bh3_w0_4 <= tile_15_filtered_output(4);
   tile_16_X <= X(5 downto 3);
   tile_16_Y <= Y(11 downto 10);
   tile_16_mult: IntMultiplierLUT_3x2_comb_uid69
      port map ( X => tile_16_X,
                 Y => tile_16_Y,
                 R => tile_16_output);

   tile_16_filtered_output <= unsigned(tile_16_output(4 downto 0));
   bh3_wm7_1 <= tile_16_filtered_output(0);
   bh3_wm6_2 <= tile_16_filtered_output(1);
   bh3_wm5_3 <= tile_16_filtered_output(2);
   bh3_wm4_4 <= tile_16_filtered_output(3);
   bh3_wm3_4 <= tile_16_filtered_output(4);
   tile_17_X <= X(2 downto 0);
   tile_17_Y <= Y(11 downto 10);
   tile_17_mult: IntMultiplierLUT_3x2_comb_uid73
      port map ( X => tile_17_X,
                 Y => tile_17_Y,
                 R => tile_17_output);

   tile_17_filtered_output <= unsigned(tile_17_output(4 downto 0));
   bh3_wm10_0 <= tile_17_filtered_output(0);
   bh3_wm9_0 <= tile_17_filtered_output(1);
   bh3_wm8_1 <= tile_17_filtered_output(2);
   bh3_wm7_2 <= tile_17_filtered_output(3);
   bh3_wm6_3 <= tile_17_filtered_output(4);
   tile_18_X <= X(15 downto 15);
   tile_18_Y <= Y(9 downto 8);
   tile_18_mult: IntMultiplierLUT_1_signedx2_comb_uid77
      port map ( X => tile_18_X,
                 Y => tile_18_Y,
                 R => tile_18_output);

   tile_18_filtered_output <= signed(tile_18_output(2 downto 0));
   bh3_w3_5 <= tile_18_filtered_output(0);
   bh3_w4_5 <= tile_18_filtered_output(1);
   bh3_w5_5 <= not tile_18_filtered_output(2);
   tile_19_X <= X(14 downto 12);
   tile_19_Y <= Y(9 downto 8);
   tile_19_mult: IntMultiplierLUT_3x2_comb_uid81
      port map ( X => tile_19_X,
                 Y => tile_19_Y,
                 R => tile_19_output);

   tile_19_filtered_output <= unsigned(tile_19_output(4 downto 0));
   bh3_w0_5 <= tile_19_filtered_output(0);
   bh3_w1_5 <= tile_19_filtered_output(1);
   bh3_w2_5 <= tile_19_filtered_output(2);
   bh3_w3_6 <= tile_19_filtered_output(3);
   bh3_w4_6 <= tile_19_filtered_output(4);
   tile_20_X <= X(11 downto 9);
   tile_20_Y <= Y(9 downto 8);
   tile_20_mult: IntMultiplierLUT_3x2_comb_uid85
      port map ( X => tile_20_X,
                 Y => tile_20_Y,
                 R => tile_20_output);

   tile_20_filtered_output <= unsigned(tile_20_output(4 downto 0));
   bh3_wm3_5 <= tile_20_filtered_output(0);
   bh3_wm2_5 <= tile_20_filtered_output(1);
   bh3_wm1_5 <= tile_20_filtered_output(2);
   bh3_w0_6 <= tile_20_filtered_output(3);
   bh3_w1_6 <= tile_20_filtered_output(4);
   tile_21_X <= X(8 downto 6);
   tile_21_Y <= Y(9 downto 8);
   tile_21_mult: IntMultiplierLUT_3x2_comb_uid89
      port map ( X => tile_21_X,
                 Y => tile_21_Y,
                 R => tile_21_output);

   tile_21_filtered_output <= unsigned(tile_21_output(4 downto 0));
   bh3_wm6_4 <= tile_21_filtered_output(0);
   bh3_wm5_4 <= tile_21_filtered_output(1);
   bh3_wm4_5 <= tile_21_filtered_output(2);
   bh3_wm3_6 <= tile_21_filtered_output(3);
   bh3_wm2_6 <= tile_21_filtered_output(4);
   tile_22_X <= X(5 downto 3);
   tile_22_Y <= Y(9 downto 8);
   tile_22_mult: IntMultiplierLUT_3x2_comb_uid93
      port map ( X => tile_22_X,
                 Y => tile_22_Y,
                 R => tile_22_output);

   tile_22_filtered_output <= unsigned(tile_22_output(4 downto 0));
   bh3_wm9_1 <= tile_22_filtered_output(0);
   bh3_wm8_2 <= tile_22_filtered_output(1);
   bh3_wm7_3 <= tile_22_filtered_output(2);
   bh3_wm6_5 <= tile_22_filtered_output(3);
   bh3_wm5_5 <= tile_22_filtered_output(4);
   tile_23_X <= X(2 downto 0);
   tile_23_Y <= Y(9 downto 8);
   tile_23_mult: IntMultiplierLUT_3x2_comb_uid97
      port map ( X => tile_23_X,
                 Y => tile_23_Y,
                 R => tile_23_output);

   tile_23_filtered_output <= unsigned(tile_23_output(4 downto 0));
   bh3_wm12_0 <= tile_23_filtered_output(0);
   bh3_wm11_0 <= tile_23_filtered_output(1);
   bh3_wm10_1 <= tile_23_filtered_output(2);
   bh3_wm9_2 <= tile_23_filtered_output(3);
   bh3_wm8_3 <= tile_23_filtered_output(4);
   tile_24_X <= X(15 downto 15);
   tile_24_Y <= Y(7 downto 6);
   tile_24_mult: IntMultiplierLUT_1_signedx2_comb_uid101
      port map ( X => tile_24_X,
                 Y => tile_24_Y,
                 R => tile_24_output);

   tile_24_filtered_output <= signed(tile_24_output(2 downto 0));
   bh3_w1_7 <= tile_24_filtered_output(0);
   bh3_w2_6 <= tile_24_filtered_output(1);
   bh3_w3_7 <= not tile_24_filtered_output(2);
   tile_25_X <= X(14 downto 12);
   tile_25_Y <= Y(7 downto 6);
   tile_25_mult: IntMultiplierLUT_3x2_comb_uid105
      port map ( X => tile_25_X,
                 Y => tile_25_Y,
                 R => tile_25_output);

   tile_25_filtered_output <= unsigned(tile_25_output(4 downto 0));
   bh3_wm2_7 <= tile_25_filtered_output(0);
   bh3_wm1_6 <= tile_25_filtered_output(1);
   bh3_w0_7 <= tile_25_filtered_output(2);
   bh3_w1_8 <= tile_25_filtered_output(3);
   bh3_w2_7 <= tile_25_filtered_output(4);
   tile_26_X <= X(11 downto 9);
   tile_26_Y <= Y(7 downto 6);
   tile_26_mult: IntMultiplierLUT_3x2_comb_uid109
      port map ( X => tile_26_X,
                 Y => tile_26_Y,
                 R => tile_26_output);

   tile_26_filtered_output <= unsigned(tile_26_output(4 downto 0));
   bh3_wm5_6 <= tile_26_filtered_output(0);
   bh3_wm4_6 <= tile_26_filtered_output(1);
   bh3_wm3_7 <= tile_26_filtered_output(2);
   bh3_wm2_8 <= tile_26_filtered_output(3);
   bh3_wm1_7 <= tile_26_filtered_output(4);
   tile_27_X <= X(8 downto 6);
   tile_27_Y <= Y(7 downto 6);
   tile_27_mult: IntMultiplierLUT_3x2_comb_uid113
      port map ( X => tile_27_X,
                 Y => tile_27_Y,
                 R => tile_27_output);

   tile_27_filtered_output <= unsigned(tile_27_output(4 downto 0));
   bh3_wm8_4 <= tile_27_filtered_output(0);
   bh3_wm7_4 <= tile_27_filtered_output(1);
   bh3_wm6_6 <= tile_27_filtered_output(2);
   bh3_wm5_7 <= tile_27_filtered_output(3);
   bh3_wm4_7 <= tile_27_filtered_output(4);
   tile_28_X <= X(5 downto 3);
   tile_28_Y <= Y(7 downto 6);
   tile_28_mult: IntMultiplierLUT_3x2_comb_uid117
      port map ( X => tile_28_X,
                 Y => tile_28_Y,
                 R => tile_28_output);

   tile_28_filtered_output <= unsigned(tile_28_output(4 downto 0));
   bh3_wm11_1 <= tile_28_filtered_output(0);
   bh3_wm10_2 <= tile_28_filtered_output(1);
   bh3_wm9_3 <= tile_28_filtered_output(2);
   bh3_wm8_5 <= tile_28_filtered_output(3);
   bh3_wm7_5 <= tile_28_filtered_output(4);
   tile_29_X <= X(2 downto 0);
   tile_29_Y <= Y(7 downto 6);
   tile_29_mult: IntMultiplierLUT_3x2_comb_uid121
      port map ( X => tile_29_X,
                 Y => tile_29_Y,
                 R => tile_29_output);

   tile_29_filtered_output <= unsigned(tile_29_output(4 downto 0));
   bh3_wm14_0 <= tile_29_filtered_output(0);
   bh3_wm13_0 <= tile_29_filtered_output(1);
   bh3_wm12_1 <= tile_29_filtered_output(2);
   bh3_wm11_2 <= tile_29_filtered_output(3);
   bh3_wm10_3 <= tile_29_filtered_output(4);
   tile_30_X <= X(15 downto 15);
   tile_30_Y <= Y(5 downto 4);
   tile_30_mult: IntMultiplierLUT_1_signedx2_comb_uid125
      port map ( X => tile_30_X,
                 Y => tile_30_Y,
                 R => tile_30_output);

   tile_30_filtered_output <= signed(tile_30_output(2 downto 0));
   bh3_wm1_8 <= tile_30_filtered_output(0);
   bh3_w0_8 <= tile_30_filtered_output(1);
   bh3_w1_9 <= not tile_30_filtered_output(2);
   tile_31_X <= X(14 downto 12);
   tile_31_Y <= Y(5 downto 4);
   tile_31_mult: IntMultiplierLUT_3x2_comb_uid129
      port map ( X => tile_31_X,
                 Y => tile_31_Y,
                 R => tile_31_output);

   tile_31_filtered_output <= unsigned(tile_31_output(4 downto 0));
   bh3_wm4_8 <= tile_31_filtered_output(0);
   bh3_wm3_8 <= tile_31_filtered_output(1);
   bh3_wm2_9 <= tile_31_filtered_output(2);
   bh3_wm1_9 <= tile_31_filtered_output(3);
   bh3_w0_9 <= tile_31_filtered_output(4);
   tile_32_X <= X(11 downto 9);
   tile_32_Y <= Y(5 downto 4);
   tile_32_mult: IntMultiplierLUT_3x2_comb_uid133
      port map ( X => tile_32_X,
                 Y => tile_32_Y,
                 R => tile_32_output);

   tile_32_filtered_output <= unsigned(tile_32_output(4 downto 0));
   bh3_wm7_6 <= tile_32_filtered_output(0);
   bh3_wm6_7 <= tile_32_filtered_output(1);
   bh3_wm5_8 <= tile_32_filtered_output(2);
   bh3_wm4_9 <= tile_32_filtered_output(3);
   bh3_wm3_9 <= tile_32_filtered_output(4);
   tile_33_X <= X(8 downto 6);
   tile_33_Y <= Y(5 downto 4);
   tile_33_mult: IntMultiplierLUT_3x2_comb_uid137
      port map ( X => tile_33_X,
                 Y => tile_33_Y,
                 R => tile_33_output);

   tile_33_filtered_output <= unsigned(tile_33_output(4 downto 0));
   bh3_wm10_4 <= tile_33_filtered_output(0);
   bh3_wm9_4 <= tile_33_filtered_output(1);
   bh3_wm8_6 <= tile_33_filtered_output(2);
   bh3_wm7_7 <= tile_33_filtered_output(3);
   bh3_wm6_8 <= tile_33_filtered_output(4);
   tile_34_X <= X(5 downto 3);
   tile_34_Y <= Y(5 downto 4);
   tile_34_mult: IntMultiplierLUT_3x2_comb_uid141
      port map ( X => tile_34_X,
                 Y => tile_34_Y,
                 R => tile_34_output);

   tile_34_filtered_output <= unsigned(tile_34_output(4 downto 0));
   bh3_wm13_1 <= tile_34_filtered_output(0);
   bh3_wm12_2 <= tile_34_filtered_output(1);
   bh3_wm11_3 <= tile_34_filtered_output(2);
   bh3_wm10_5 <= tile_34_filtered_output(3);
   bh3_wm9_5 <= tile_34_filtered_output(4);
   tile_35_X <= X(2 downto 0);
   tile_35_Y <= Y(5 downto 4);
   tile_35_mult: IntMultiplierLUT_3x2_comb_uid145
      port map ( X => tile_35_X,
                 Y => tile_35_Y,
                 R => tile_35_output);

   tile_35_filtered_output <= unsigned(tile_35_output(4 downto 0));
   bh3_wm16_0 <= tile_35_filtered_output(0);
   bh3_wm15_0 <= tile_35_filtered_output(1);
   bh3_wm14_1 <= tile_35_filtered_output(2);
   bh3_wm13_2 <= tile_35_filtered_output(3);
   bh3_wm12_3 <= tile_35_filtered_output(4);
   tile_36_X <= X(15 downto 15);
   tile_36_Y <= Y(3 downto 2);
   tile_36_mult: IntMultiplierLUT_1_signedx2_comb_uid149
      port map ( X => tile_36_X,
                 Y => tile_36_Y,
                 R => tile_36_output);

   tile_36_filtered_output <= signed(tile_36_output(2 downto 0));
   bh3_wm3_10 <= tile_36_filtered_output(0);
   bh3_wm2_10 <= tile_36_filtered_output(1);
   bh3_wm1_10 <= not tile_36_filtered_output(2);
   tile_37_X <= X(14 downto 12);
   tile_37_Y <= Y(3 downto 2);
   tile_37_mult: IntMultiplierLUT_3x2_comb_uid153
      port map ( X => tile_37_X,
                 Y => tile_37_Y,
                 R => tile_37_output);

   tile_37_filtered_output <= unsigned(tile_37_output(4 downto 0));
   bh3_wm6_9 <= tile_37_filtered_output(0);
   bh3_wm5_9 <= tile_37_filtered_output(1);
   bh3_wm4_10 <= tile_37_filtered_output(2);
   bh3_wm3_11 <= tile_37_filtered_output(3);
   bh3_wm2_11 <= tile_37_filtered_output(4);
   tile_38_X <= X(11 downto 9);
   tile_38_Y <= Y(3 downto 2);
   tile_38_mult: IntMultiplierLUT_3x2_comb_uid157
      port map ( X => tile_38_X,
                 Y => tile_38_Y,
                 R => tile_38_output);

   tile_38_filtered_output <= unsigned(tile_38_output(4 downto 0));
   bh3_wm9_6 <= tile_38_filtered_output(0);
   bh3_wm8_7 <= tile_38_filtered_output(1);
   bh3_wm7_8 <= tile_38_filtered_output(2);
   bh3_wm6_10 <= tile_38_filtered_output(3);
   bh3_wm5_10 <= tile_38_filtered_output(4);
   tile_39_X <= X(8 downto 6);
   tile_39_Y <= Y(3 downto 2);
   tile_39_mult: IntMultiplierLUT_3x2_comb_uid161
      port map ( X => tile_39_X,
                 Y => tile_39_Y,
                 R => tile_39_output);

   tile_39_filtered_output <= unsigned(tile_39_output(4 downto 0));
   bh3_wm12_4 <= tile_39_filtered_output(0);
   bh3_wm11_4 <= tile_39_filtered_output(1);
   bh3_wm10_6 <= tile_39_filtered_output(2);
   bh3_wm9_7 <= tile_39_filtered_output(3);
   bh3_wm8_8 <= tile_39_filtered_output(4);
   tile_40_X <= X(5 downto 3);
   tile_40_Y <= Y(3 downto 2);
   tile_40_mult: IntMultiplierLUT_3x2_comb_uid165
      port map ( X => tile_40_X,
                 Y => tile_40_Y,
                 R => tile_40_output);

   tile_40_filtered_output <= unsigned(tile_40_output(4 downto 0));
   bh3_wm15_1 <= tile_40_filtered_output(0);
   bh3_wm14_2 <= tile_40_filtered_output(1);
   bh3_wm13_3 <= tile_40_filtered_output(2);
   bh3_wm12_5 <= tile_40_filtered_output(3);
   bh3_wm11_5 <= tile_40_filtered_output(4);
   tile_41_X <= X(2 downto 0);
   tile_41_Y <= Y(3 downto 2);
   tile_41_mult: IntMultiplierLUT_3x2_comb_uid169
      port map ( X => tile_41_X,
                 Y => tile_41_Y,
                 R => tile_41_output);

   tile_41_filtered_output <= unsigned(tile_41_output(4 downto 0));
   bh3_wm18_0 <= tile_41_filtered_output(0);
   bh3_wm17_0 <= tile_41_filtered_output(1);
   bh3_wm16_1 <= tile_41_filtered_output(2);
   bh3_wm15_2 <= tile_41_filtered_output(3);
   bh3_wm14_3 <= tile_41_filtered_output(4);
   tile_42_X <= X(15 downto 15);
   tile_42_Y <= Y(1 downto 0);
   tile_42_mult: IntMultiplierLUT_1_signedx2_comb_uid173
      port map ( X => tile_42_X,
                 Y => tile_42_Y,
                 R => tile_42_output);

   tile_42_filtered_output <= signed(tile_42_output(2 downto 0));
   bh3_wm5_11 <= tile_42_filtered_output(0);
   bh3_wm4_11 <= tile_42_filtered_output(1);
   bh3_wm3_12 <= not tile_42_filtered_output(2);
   tile_43_X <= X(14 downto 12);
   tile_43_Y <= Y(1 downto 0);
   tile_43_mult: IntMultiplierLUT_3x2_comb_uid177
      port map ( X => tile_43_X,
                 Y => tile_43_Y,
                 R => tile_43_output);

   tile_43_filtered_output <= unsigned(tile_43_output(4 downto 0));
   bh3_wm8_9 <= tile_43_filtered_output(0);
   bh3_wm7_9 <= tile_43_filtered_output(1);
   bh3_wm6_11 <= tile_43_filtered_output(2);
   bh3_wm5_12 <= tile_43_filtered_output(3);
   bh3_wm4_12 <= tile_43_filtered_output(4);
   tile_44_X <= X(11 downto 9);
   tile_44_Y <= Y(1 downto 0);
   tile_44_mult: IntMultiplierLUT_3x2_comb_uid181
      port map ( X => tile_44_X,
                 Y => tile_44_Y,
                 R => tile_44_output);

   tile_44_filtered_output <= unsigned(tile_44_output(4 downto 0));
   bh3_wm11_6 <= tile_44_filtered_output(0);
   bh3_wm10_7 <= tile_44_filtered_output(1);
   bh3_wm9_8 <= tile_44_filtered_output(2);
   bh3_wm8_10 <= tile_44_filtered_output(3);
   bh3_wm7_10 <= tile_44_filtered_output(4);
   tile_45_X <= X(8 downto 6);
   tile_45_Y <= Y(1 downto 0);
   tile_45_mult: IntMultiplierLUT_3x2_comb_uid185
      port map ( X => tile_45_X,
                 Y => tile_45_Y,
                 R => tile_45_output);

   tile_45_filtered_output <= unsigned(tile_45_output(4 downto 0));
   bh3_wm14_4 <= tile_45_filtered_output(0);
   bh3_wm13_4 <= tile_45_filtered_output(1);
   bh3_wm12_6 <= tile_45_filtered_output(2);
   bh3_wm11_7 <= tile_45_filtered_output(3);
   bh3_wm10_8 <= tile_45_filtered_output(4);
   tile_46_X <= X(5 downto 3);
   tile_46_Y <= Y(1 downto 0);
   tile_46_mult: IntMultiplierLUT_3x2_comb_uid189
      port map ( X => tile_46_X,
                 Y => tile_46_Y,
                 R => tile_46_output);

   tile_46_filtered_output <= unsigned(tile_46_output(4 downto 0));
   bh3_wm17_1 <= tile_46_filtered_output(0);
   bh3_wm16_2 <= tile_46_filtered_output(1);
   bh3_wm15_3 <= tile_46_filtered_output(2);
   bh3_wm14_5 <= tile_46_filtered_output(3);
   bh3_wm13_5 <= tile_46_filtered_output(4);
   tile_47_X <= X(2 downto 0);
   tile_47_Y <= Y(1 downto 0);
   tile_47_mult: IntMultiplierLUT_3x2_comb_uid193
      port map ( X => tile_47_X,
                 Y => tile_47_Y,
                 R => tile_47_output);

   tile_47_filtered_output <= unsigned(tile_47_output(4 downto 0));
   bh3_wm20_0 <= tile_47_filtered_output(0);
   bh3_wm19_0 <= tile_47_filtered_output(1);
   bh3_wm18_1 <= tile_47_filtered_output(2);
   bh3_wm17_2 <= tile_47_filtered_output(3);
   bh3_wm16_3 <= tile_47_filtered_output(4);
   bh3_wm20_1 <= AA(0);
   bh3_wm19_1 <= AA(1);
   bh3_wm18_2 <= AA(2);
   bh3_wm17_3 <= AA(3);
   bh3_wm16_4 <= AA(4);
   bh3_wm15_4 <= AA(5);
   bh3_wm14_6 <= AA(6);
   bh3_wm13_6 <= AA(7);
   bh3_wm12_7 <= AA(8);
   bh3_wm11_8 <= AA(9);
   bh3_wm10_9 <= AA(10);
   bh3_wm9_9 <= AA(11);
   bh3_wm8_11 <= AA(12);
   bh3_wm7_11 <= AA(13);
   bh3_wm6_12 <= AA(14);
   bh3_wm5_13 <= AA(15);
   bh3_wm4_13 <= AA(16);
   bh3_wm3_13 <= AA(17);
   bh3_wm2_12 <= AA(18);
   bh3_wm1_11 <= AA(19);
   bh3_w0_10 <= AA(20);
   bh3_w1_10 <= AA(21);
   bh3_w2_8 <= AA(22);
   bh3_w3_8 <= AA(23);
   bh3_w4_7 <= AA(24);
   bh3_w5_6 <= AA(25);
   bh3_w6_5 <= AA(26);
   bh3_w7_5 <= AA(27);
   bh3_w8_3 <= AA(28);
   bh3_w9_3 <= AA(29);
   bh3_w10_2 <= AA(30);
   bh3_w11_1 <= AA(31);

   -- Adding the constant bits 
   bh3_wm3_14 <= '1';
   bh3_w0_11 <= '1';
   bh3_w1_11 <= '1';
   bh3_w6_6 <= '1';
   bh3_w7_6 <= '1';


   Compressor_23_3_comb_uid198_bh3_uid199_In0 <= "" & bh3_wm20_1 & bh3_wm20_0 & "0";
   Compressor_23_3_comb_uid198_bh3_uid199_In1 <= "" & bh3_wm19_1 & bh3_wm19_0;
   bh3_wm20_2 <= Compressor_23_3_comb_uid198_bh3_uid199_Out0(0);
   bh3_wm19_2 <= Compressor_23_3_comb_uid198_bh3_uid199_Out0(1);
   bh3_wm18_3 <= Compressor_23_3_comb_uid198_bh3_uid199_Out0(2);
   Compressor_23_3_comb_uid198_uid199: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid199_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid199_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid199_Out0);


   Compressor_3_2_comb_uid201_bh3_uid202_In0 <= "" & bh3_wm18_2 & bh3_wm18_0 & bh3_wm18_1;
   bh3_wm18_4 <= Compressor_3_2_comb_uid201_bh3_uid202_Out0(0);
   bh3_wm17_4 <= Compressor_3_2_comb_uid201_bh3_uid202_Out0(1);
   Compressor_3_2_comb_uid201_uid202: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid202_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid202_Out0);


   Compressor_14_3_comb_uid204_bh3_uid205_In0 <= "" & bh3_wm17_3 & bh3_wm17_0 & bh3_wm17_1 & bh3_wm17_2;
   Compressor_14_3_comb_uid204_bh3_uid205_In1 <= "" & bh3_wm16_4;
   bh3_wm17_5 <= Compressor_14_3_comb_uid204_bh3_uid205_Out0(0);
   bh3_wm16_5 <= Compressor_14_3_comb_uid204_bh3_uid205_Out0(1);
   bh3_wm15_5 <= Compressor_14_3_comb_uid204_bh3_uid205_Out0(2);
   Compressor_14_3_comb_uid204_uid205: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid205_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid205_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid205_Out0);


   Compressor_14_3_comb_uid204_bh3_uid206_In0 <= "" & bh3_wm16_0 & bh3_wm16_1 & bh3_wm16_2 & bh3_wm16_3;
   Compressor_14_3_comb_uid204_bh3_uid206_In1 <= "" & bh3_wm15_4;
   bh3_wm16_6 <= Compressor_14_3_comb_uid204_bh3_uid206_Out0(0);
   bh3_wm15_6 <= Compressor_14_3_comb_uid204_bh3_uid206_Out0(1);
   bh3_wm14_7 <= Compressor_14_3_comb_uid204_bh3_uid206_Out0(2);
   Compressor_14_3_comb_uid204_uid206: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid206_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid206_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid206_Out0);


   Compressor_14_3_comb_uid204_bh3_uid207_In0 <= "" & bh3_wm15_0 & bh3_wm15_1 & bh3_wm15_2 & bh3_wm15_3;
   Compressor_14_3_comb_uid204_bh3_uid207_In1 <= "" & bh3_wm14_6;
   bh3_wm15_7 <= Compressor_14_3_comb_uid204_bh3_uid207_Out0(0);
   bh3_wm14_8 <= Compressor_14_3_comb_uid204_bh3_uid207_Out0(1);
   bh3_wm13_7 <= Compressor_14_3_comb_uid204_bh3_uid207_Out0(2);
   Compressor_14_3_comb_uid204_uid207: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid207_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid207_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid207_Out0);


   Compressor_6_3_comb_uid209_bh3_uid210_In0 <= "" & bh3_wm14_0 & bh3_wm14_1 & bh3_wm14_2 & bh3_wm14_3 & bh3_wm14_4 & bh3_wm14_5;
   bh3_wm14_9 <= Compressor_6_3_comb_uid209_bh3_uid210_Out0(0);
   bh3_wm13_8 <= Compressor_6_3_comb_uid209_bh3_uid210_Out0(1);
   bh3_wm12_8 <= Compressor_6_3_comb_uid209_bh3_uid210_Out0(2);
   Compressor_6_3_comb_uid209_uid210: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid210_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid210_Out0);


   Compressor_6_3_comb_uid209_bh3_uid211_In0 <= "" & bh3_wm13_6 & bh3_wm13_0 & bh3_wm13_1 & bh3_wm13_2 & "0" & "0";
   bh3_wm13_9 <= Compressor_6_3_comb_uid209_bh3_uid211_Out0(0);
   bh3_wm12_9 <= Compressor_6_3_comb_uid209_bh3_uid211_Out0(1);
   bh3_wm11_9 <= Compressor_6_3_comb_uid209_bh3_uid211_Out0(2);
   Compressor_6_3_comb_uid209_uid211: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid211_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid211_Out0);


   Compressor_23_3_comb_uid198_bh3_uid212_In0 <= "" & bh3_wm13_3 & bh3_wm13_4 & bh3_wm13_5;
   Compressor_23_3_comb_uid198_bh3_uid212_In1 <= "" & bh3_wm12_7 & bh3_wm12_0;
   bh3_wm13_10 <= Compressor_23_3_comb_uid198_bh3_uid212_Out0(0);
   bh3_wm12_10 <= Compressor_23_3_comb_uid198_bh3_uid212_Out0(1);
   bh3_wm11_10 <= Compressor_23_3_comb_uid198_bh3_uid212_Out0(2);
   Compressor_23_3_comb_uid198_uid212: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid212_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid212_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid212_Out0);


   Compressor_6_3_comb_uid209_bh3_uid213_In0 <= "" & bh3_wm12_1 & bh3_wm12_2 & bh3_wm12_3 & bh3_wm12_4 & bh3_wm12_5 & bh3_wm12_6;
   bh3_wm12_11 <= Compressor_6_3_comb_uid209_bh3_uid213_Out0(0);
   bh3_wm11_11 <= Compressor_6_3_comb_uid209_bh3_uid213_Out0(1);
   bh3_wm10_10 <= Compressor_6_3_comb_uid209_bh3_uid213_Out0(2);
   Compressor_6_3_comb_uid209_uid213: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid213_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid213_Out0);


   Compressor_6_3_comb_uid209_bh3_uid214_In0 <= "" & bh3_wm11_8 & bh3_wm11_0 & bh3_wm11_1 & bh3_wm11_2 & bh3_wm11_3 & bh3_wm11_4;
   bh3_wm11_12 <= Compressor_6_3_comb_uid209_bh3_uid214_Out0(0);
   bh3_wm10_11 <= Compressor_6_3_comb_uid209_bh3_uid214_Out0(1);
   bh3_wm9_10 <= Compressor_6_3_comb_uid209_bh3_uid214_Out0(2);
   Compressor_6_3_comb_uid209_uid214: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid214_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid214_Out0);


   Compressor_3_2_comb_uid201_bh3_uid215_In0 <= "" & bh3_wm11_5 & bh3_wm11_6 & bh3_wm11_7;
   bh3_wm11_13 <= Compressor_3_2_comb_uid201_bh3_uid215_Out0(0);
   bh3_wm10_12 <= Compressor_3_2_comb_uid201_bh3_uid215_Out0(1);
   Compressor_3_2_comb_uid201_uid215: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid215_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid215_Out0);


   Compressor_6_3_comb_uid209_bh3_uid216_In0 <= "" & bh3_wm10_9 & bh3_wm10_0 & bh3_wm10_1 & bh3_wm10_2 & bh3_wm10_3 & bh3_wm10_4;
   bh3_wm10_13 <= Compressor_6_3_comb_uid209_bh3_uid216_Out0(0);
   bh3_wm9_11 <= Compressor_6_3_comb_uid209_bh3_uid216_Out0(1);
   bh3_wm8_12 <= Compressor_6_3_comb_uid209_bh3_uid216_Out0(2);
   Compressor_6_3_comb_uid209_uid216: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid216_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid216_Out0);


   Compressor_14_3_comb_uid204_bh3_uid217_In0 <= "" & bh3_wm10_5 & bh3_wm10_6 & bh3_wm10_7 & bh3_wm10_8;
   Compressor_14_3_comb_uid204_bh3_uid217_In1 <= "" & bh3_wm9_9;
   bh3_wm10_14 <= Compressor_14_3_comb_uid204_bh3_uid217_Out0(0);
   bh3_wm9_12 <= Compressor_14_3_comb_uid204_bh3_uid217_Out0(1);
   bh3_wm8_13 <= Compressor_14_3_comb_uid204_bh3_uid217_Out0(2);
   Compressor_14_3_comb_uid204_uid217: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid217_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid217_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid217_Out0);


   Compressor_6_3_comb_uid209_bh3_uid218_In0 <= "" & bh3_wm9_0 & bh3_wm9_1 & bh3_wm9_2 & bh3_wm9_3 & bh3_wm9_4 & bh3_wm9_5;
   bh3_wm9_13 <= Compressor_6_3_comb_uid209_bh3_uid218_Out0(0);
   bh3_wm8_14 <= Compressor_6_3_comb_uid209_bh3_uid218_Out0(1);
   bh3_wm7_12 <= Compressor_6_3_comb_uid209_bh3_uid218_Out0(2);
   Compressor_6_3_comb_uid209_uid218: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid218_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid218_Out0);


   Compressor_3_2_comb_uid201_bh3_uid219_In0 <= "" & bh3_wm9_6 & bh3_wm9_7 & bh3_wm9_8;
   bh3_wm9_14 <= Compressor_3_2_comb_uid201_bh3_uid219_Out0(0);
   bh3_wm8_15 <= Compressor_3_2_comb_uid201_bh3_uid219_Out0(1);
   Compressor_3_2_comb_uid201_uid219: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid219_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid219_Out0);


   Compressor_6_3_comb_uid209_bh3_uid220_In0 <= "" & bh3_wm8_11 & bh3_wm8_0 & bh3_wm8_1 & bh3_wm8_2 & bh3_wm8_3 & bh3_wm8_4;
   bh3_wm8_16 <= Compressor_6_3_comb_uid209_bh3_uid220_Out0(0);
   bh3_wm7_13 <= Compressor_6_3_comb_uid209_bh3_uid220_Out0(1);
   bh3_wm6_13 <= Compressor_6_3_comb_uid209_bh3_uid220_Out0(2);
   Compressor_6_3_comb_uid209_uid220: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid220_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid220_Out0);


   Compressor_6_3_comb_uid209_bh3_uid221_In0 <= "" & bh3_wm8_5 & bh3_wm8_6 & bh3_wm8_7 & bh3_wm8_8 & bh3_wm8_9 & bh3_wm8_10;
   bh3_wm8_17 <= Compressor_6_3_comb_uid209_bh3_uid221_Out0(0);
   bh3_wm7_14 <= Compressor_6_3_comb_uid209_bh3_uid221_Out0(1);
   bh3_wm6_14 <= Compressor_6_3_comb_uid209_bh3_uid221_Out0(2);
   Compressor_6_3_comb_uid209_uid221: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid221_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid221_Out0);


   Compressor_6_3_comb_uid209_bh3_uid222_In0 <= "" & bh3_wm7_11 & bh3_wm7_0 & bh3_wm7_1 & bh3_wm7_2 & bh3_wm7_3 & bh3_wm7_4;
   bh3_wm7_15 <= Compressor_6_3_comb_uid209_bh3_uid222_Out0(0);
   bh3_wm6_15 <= Compressor_6_3_comb_uid209_bh3_uid222_Out0(1);
   bh3_wm5_14 <= Compressor_6_3_comb_uid209_bh3_uid222_Out0(2);
   Compressor_6_3_comb_uid209_uid222: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid222_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid222_Out0);


   Compressor_6_3_comb_uid209_bh3_uid223_In0 <= "" & bh3_wm7_5 & bh3_wm7_6 & bh3_wm7_7 & bh3_wm7_8 & bh3_wm7_9 & bh3_wm7_10;
   bh3_wm7_16 <= Compressor_6_3_comb_uid209_bh3_uid223_Out0(0);
   bh3_wm6_16 <= Compressor_6_3_comb_uid209_bh3_uid223_Out0(1);
   bh3_wm5_15 <= Compressor_6_3_comb_uid209_bh3_uid223_Out0(2);
   Compressor_6_3_comb_uid209_uid223: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid223_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid223_Out0);


   Compressor_6_3_comb_uid209_bh3_uid224_In0 <= "" & bh3_wm6_12 & bh3_wm6_0 & bh3_wm6_1 & bh3_wm6_2 & bh3_wm6_3 & bh3_wm6_4;
   bh3_wm6_17 <= Compressor_6_3_comb_uid209_bh3_uid224_Out0(0);
   bh3_wm5_16 <= Compressor_6_3_comb_uid209_bh3_uid224_Out0(1);
   bh3_wm4_14 <= Compressor_6_3_comb_uid209_bh3_uid224_Out0(2);
   Compressor_6_3_comb_uid209_uid224: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid224_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid224_Out0);


   Compressor_6_3_comb_uid209_bh3_uid225_In0 <= "" & bh3_wm6_5 & bh3_wm6_6 & bh3_wm6_7 & bh3_wm6_8 & bh3_wm6_9 & bh3_wm6_10;
   bh3_wm6_18 <= Compressor_6_3_comb_uid209_bh3_uid225_Out0(0);
   bh3_wm5_17 <= Compressor_6_3_comb_uid209_bh3_uid225_Out0(1);
   bh3_wm4_15 <= Compressor_6_3_comb_uid209_bh3_uid225_Out0(2);
   Compressor_6_3_comb_uid209_uid225: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid225_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid225_Out0);


   Compressor_6_3_comb_uid209_bh3_uid226_In0 <= "" & bh3_wm5_13 & bh3_wm5_0 & bh3_wm5_1 & bh3_wm5_2 & bh3_wm5_3 & "0";
   bh3_wm5_18 <= Compressor_6_3_comb_uid209_bh3_uid226_Out0(0);
   bh3_wm4_16 <= Compressor_6_3_comb_uid209_bh3_uid226_Out0(1);
   bh3_wm3_15 <= Compressor_6_3_comb_uid209_bh3_uid226_Out0(2);
   Compressor_6_3_comb_uid209_uid226: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid226_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid226_Out0);


   Compressor_6_3_comb_uid209_bh3_uid227_In0 <= "" & bh3_wm5_4 & bh3_wm5_5 & bh3_wm5_6 & bh3_wm5_7 & bh3_wm5_8 & bh3_wm5_9;
   bh3_wm5_19 <= Compressor_6_3_comb_uid209_bh3_uid227_Out0(0);
   bh3_wm4_17 <= Compressor_6_3_comb_uid209_bh3_uid227_Out0(1);
   bh3_wm3_16 <= Compressor_6_3_comb_uid209_bh3_uid227_Out0(2);
   Compressor_6_3_comb_uid209_uid227: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid227_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid227_Out0);


   Compressor_23_3_comb_uid198_bh3_uid228_In0 <= "" & bh3_wm5_12 & bh3_wm5_11 & bh3_wm5_10;
   Compressor_23_3_comb_uid198_bh3_uid228_In1 <= "" & bh3_wm4_13 & bh3_wm4_0;
   bh3_wm5_20 <= Compressor_23_3_comb_uid198_bh3_uid228_Out0(0);
   bh3_wm4_18 <= Compressor_23_3_comb_uid198_bh3_uid228_Out0(1);
   bh3_wm3_17 <= Compressor_23_3_comb_uid198_bh3_uid228_Out0(2);
   Compressor_23_3_comb_uid198_uid228: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid228_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid228_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid228_Out0);


   Compressor_6_3_comb_uid209_bh3_uid229_In0 <= "" & bh3_wm4_1 & bh3_wm4_2 & bh3_wm4_3 & bh3_wm4_4 & bh3_wm4_5 & bh3_wm4_6;
   bh3_wm4_19 <= Compressor_6_3_comb_uid209_bh3_uid229_Out0(0);
   bh3_wm3_18 <= Compressor_6_3_comb_uid209_bh3_uid229_Out0(1);
   bh3_wm2_13 <= Compressor_6_3_comb_uid209_bh3_uid229_Out0(2);
   Compressor_6_3_comb_uid209_uid229: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid229_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid229_Out0);


   Compressor_6_3_comb_uid209_bh3_uid230_In0 <= "" & bh3_wm4_12 & bh3_wm4_11 & bh3_wm4_10 & bh3_wm4_9 & bh3_wm4_8 & bh3_wm4_7;
   bh3_wm4_20 <= Compressor_6_3_comb_uid209_bh3_uid230_Out0(0);
   bh3_wm3_19 <= Compressor_6_3_comb_uid209_bh3_uid230_Out0(1);
   bh3_wm2_14 <= Compressor_6_3_comb_uid209_bh3_uid230_Out0(2);
   Compressor_6_3_comb_uid209_uid230: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid230_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid230_Out0);


   Compressor_6_3_comb_uid209_bh3_uid231_In0 <= "" & bh3_wm3_13 & bh3_wm3_14 & bh3_wm3_4 & bh3_wm3_7 & bh3_wm3_0 & bh3_wm3_1;
   bh3_wm3_20 <= Compressor_6_3_comb_uid209_bh3_uid231_Out0(0);
   bh3_wm2_15 <= Compressor_6_3_comb_uid209_bh3_uid231_Out0(1);
   bh3_wm1_12 <= Compressor_6_3_comb_uid209_bh3_uid231_Out0(2);
   Compressor_6_3_comb_uid209_uid231: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid231_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid231_Out0);


   Compressor_6_3_comb_uid209_bh3_uid232_In0 <= "" & bh3_wm3_9 & bh3_wm3_6 & bh3_wm3_5 & bh3_wm3_12 & bh3_wm3_11 & bh3_wm3_10;
   bh3_wm3_21 <= Compressor_6_3_comb_uid209_bh3_uid232_Out0(0);
   bh3_wm2_16 <= Compressor_6_3_comb_uid209_bh3_uid232_Out0(1);
   bh3_wm1_13 <= Compressor_6_3_comb_uid209_bh3_uid232_Out0(2);
   Compressor_6_3_comb_uid209_uid232: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid232_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid232_Out0);


   Compressor_3_2_comb_uid201_bh3_uid233_In0 <= "" & bh3_wm3_2 & bh3_wm3_3 & bh3_wm3_8;
   bh3_wm3_22 <= Compressor_3_2_comb_uid201_bh3_uid233_Out0(0);
   bh3_wm2_17 <= Compressor_3_2_comb_uid201_bh3_uid233_Out0(1);
   Compressor_3_2_comb_uid201_uid233: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid233_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid233_Out0);


   Compressor_6_3_comb_uid209_bh3_uid234_In0 <= "" & bh3_wm2_12 & bh3_wm2_0 & bh3_wm2_1 & bh3_wm2_2 & bh3_wm2_3 & bh3_wm2_4;
   bh3_wm2_18 <= Compressor_6_3_comb_uid209_bh3_uid234_Out0(0);
   bh3_wm1_14 <= Compressor_6_3_comb_uid209_bh3_uid234_Out0(1);
   bh3_w0_12 <= Compressor_6_3_comb_uid209_bh3_uid234_Out0(2);
   Compressor_6_3_comb_uid209_uid234: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid234_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid234_Out0);


   Compressor_6_3_comb_uid209_bh3_uid235_In0 <= "" & bh3_wm2_5 & bh3_wm2_6 & bh3_wm2_7 & bh3_wm2_8 & bh3_wm2_9 & bh3_wm2_10;
   bh3_wm2_19 <= Compressor_6_3_comb_uid209_bh3_uid235_Out0(0);
   bh3_wm1_15 <= Compressor_6_3_comb_uid209_bh3_uid235_Out0(1);
   bh3_w0_13 <= Compressor_6_3_comb_uid209_bh3_uid235_Out0(2);
   Compressor_6_3_comb_uid209_uid235: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid235_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid235_Out0);


   Compressor_6_3_comb_uid209_bh3_uid236_In0 <= "" & bh3_wm1_11 & bh3_wm1_0 & bh3_wm1_1 & bh3_wm1_2 & bh3_wm1_3 & bh3_wm1_4;
   bh3_wm1_16 <= Compressor_6_3_comb_uid209_bh3_uid236_Out0(0);
   bh3_w0_14 <= Compressor_6_3_comb_uid209_bh3_uid236_Out0(1);
   bh3_w1_12 <= Compressor_6_3_comb_uid209_bh3_uid236_Out0(2);
   Compressor_6_3_comb_uid209_uid236: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid236_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid236_Out0);


   Compressor_6_3_comb_uid209_bh3_uid237_In0 <= "" & bh3_wm1_5 & bh3_wm1_6 & bh3_wm1_7 & bh3_wm1_8 & bh3_wm1_9 & bh3_wm1_10;
   bh3_wm1_17 <= Compressor_6_3_comb_uid209_bh3_uid237_Out0(0);
   bh3_w0_15 <= Compressor_6_3_comb_uid209_bh3_uid237_Out0(1);
   bh3_w1_13 <= Compressor_6_3_comb_uid209_bh3_uid237_Out0(2);
   Compressor_6_3_comb_uid209_uid237: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid237_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid237_Out0);


   Compressor_6_3_comb_uid209_bh3_uid238_In0 <= "" & bh3_w0_10 & bh3_w0_11 & bh3_w0_0 & bh3_w0_1 & bh3_w0_2 & bh3_w0_3;
   bh3_w0_16 <= Compressor_6_3_comb_uid209_bh3_uid238_Out0(0);
   bh3_w1_14 <= Compressor_6_3_comb_uid209_bh3_uid238_Out0(1);
   bh3_w2_9 <= Compressor_6_3_comb_uid209_bh3_uid238_Out0(2);
   Compressor_6_3_comb_uid209_uid238: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid238_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid238_Out0);


   Compressor_6_3_comb_uid209_bh3_uid239_In0 <= "" & bh3_w0_5 & bh3_w0_9 & bh3_w0_8 & bh3_w0_7 & bh3_w0_6 & bh3_w0_4;
   bh3_w0_17 <= Compressor_6_3_comb_uid209_bh3_uid239_Out0(0);
   bh3_w1_15 <= Compressor_6_3_comb_uid209_bh3_uid239_Out0(1);
   bh3_w2_10 <= Compressor_6_3_comb_uid209_bh3_uid239_Out0(2);
   Compressor_6_3_comb_uid209_uid239: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid239_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid239_Out0);


   Compressor_6_3_comb_uid209_bh3_uid240_In0 <= "" & bh3_w1_10 & bh3_w1_11 & bh3_w1_0 & bh3_w1_1 & bh3_w1_2 & bh3_w1_3;
   bh3_w1_16 <= Compressor_6_3_comb_uid209_bh3_uid240_Out0(0);
   bh3_w2_11 <= Compressor_6_3_comb_uid209_bh3_uid240_Out0(1);
   bh3_w3_9 <= Compressor_6_3_comb_uid209_bh3_uid240_Out0(2);
   Compressor_6_3_comb_uid209_uid240: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid240_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid240_Out0);


   Compressor_6_3_comb_uid209_bh3_uid241_In0 <= "" & bh3_w1_5 & bh3_w1_9 & bh3_w1_8 & bh3_w1_7 & bh3_w1_6 & bh3_w1_4;
   bh3_w1_17 <= Compressor_6_3_comb_uid209_bh3_uid241_Out0(0);
   bh3_w2_12 <= Compressor_6_3_comb_uid209_bh3_uid241_Out0(1);
   bh3_w3_10 <= Compressor_6_3_comb_uid209_bh3_uid241_Out0(2);
   Compressor_6_3_comb_uid209_uid241: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid241_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid241_Out0);


   Compressor_6_3_comb_uid209_bh3_uid242_In0 <= "" & bh3_w2_8 & bh3_w2_0 & bh3_w2_1 & bh3_w2_2 & bh3_w2_3 & bh3_w2_4;
   bh3_w2_13 <= Compressor_6_3_comb_uid209_bh3_uid242_Out0(0);
   bh3_w3_11 <= Compressor_6_3_comb_uid209_bh3_uid242_Out0(1);
   bh3_w4_8 <= Compressor_6_3_comb_uid209_bh3_uid242_Out0(2);
   Compressor_6_3_comb_uid209_uid242: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid242_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid242_Out0);


   Compressor_23_3_comb_uid198_bh3_uid243_In0 <= "" & bh3_w2_5 & bh3_w2_6 & bh3_w2_7;
   Compressor_23_3_comb_uid198_bh3_uid243_In1 <= "" & bh3_w3_8 & bh3_w3_0;
   bh3_w2_14 <= Compressor_23_3_comb_uid198_bh3_uid243_Out0(0);
   bh3_w3_12 <= Compressor_23_3_comb_uid198_bh3_uid243_Out0(1);
   bh3_w4_9 <= Compressor_23_3_comb_uid198_bh3_uid243_Out0(2);
   Compressor_23_3_comb_uid198_uid243: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid243_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid243_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid243_Out0);


   Compressor_6_3_comb_uid209_bh3_uid244_In0 <= "" & bh3_w3_1 & bh3_w3_2 & bh3_w3_3 & bh3_w3_4 & bh3_w3_5 & bh3_w3_6;
   bh3_w3_13 <= Compressor_6_3_comb_uid209_bh3_uid244_Out0(0);
   bh3_w4_10 <= Compressor_6_3_comb_uid209_bh3_uid244_Out0(1);
   bh3_w5_7 <= Compressor_6_3_comb_uid209_bh3_uid244_Out0(2);
   Compressor_6_3_comb_uid209_uid244: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid244_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid244_Out0);


   Compressor_6_3_comb_uid209_bh3_uid245_In0 <= "" & bh3_w4_7 & bh3_w4_0 & bh3_w4_1 & bh3_w4_2 & "0" & "0";
   bh3_w4_11 <= Compressor_6_3_comb_uid209_bh3_uid245_Out0(0);
   bh3_w5_8 <= Compressor_6_3_comb_uid209_bh3_uid245_Out0(1);
   bh3_w6_7 <= Compressor_6_3_comb_uid209_bh3_uid245_Out0(2);
   Compressor_6_3_comb_uid209_uid245: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid245_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid245_Out0);


   Compressor_14_3_comb_uid204_bh3_uid246_In0 <= "" & bh3_w4_3 & bh3_w4_4 & bh3_w4_5 & bh3_w4_6;
   Compressor_14_3_comb_uid204_bh3_uid246_In1 <= "" & bh3_w5_6;
   bh3_w4_12 <= Compressor_14_3_comb_uid204_bh3_uid246_Out0(0);
   bh3_w5_9 <= Compressor_14_3_comb_uid204_bh3_uid246_Out0(1);
   bh3_w6_8 <= Compressor_14_3_comb_uid204_bh3_uid246_Out0(2);
   Compressor_14_3_comb_uid204_uid246: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid246_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid246_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid246_Out0);


   Compressor_6_3_comb_uid209_bh3_uid247_In0 <= "" & bh3_w5_0 & bh3_w5_1 & bh3_w5_2 & bh3_w5_3 & bh3_w5_4 & bh3_w5_5;
   bh3_w5_10 <= Compressor_6_3_comb_uid209_bh3_uid247_Out0(0);
   bh3_w6_9 <= Compressor_6_3_comb_uid209_bh3_uid247_Out0(1);
   bh3_w7_7 <= Compressor_6_3_comb_uid209_bh3_uid247_Out0(2);
   Compressor_6_3_comb_uid209_uid247: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid247_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid247_Out0);


   Compressor_6_3_comb_uid209_bh3_uid248_In0 <= "" & bh3_w6_5 & bh3_w6_6 & bh3_w6_0 & bh3_w6_1 & bh3_w6_2 & bh3_w6_3;
   bh3_w6_10 <= Compressor_6_3_comb_uid209_bh3_uid248_Out0(0);
   bh3_w7_8 <= Compressor_6_3_comb_uid209_bh3_uid248_Out0(1);
   bh3_w8_4 <= Compressor_6_3_comb_uid209_bh3_uid248_Out0(2);
   Compressor_6_3_comb_uid209_uid248: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid248_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid248_Out0);


   Compressor_6_3_comb_uid209_bh3_uid249_In0 <= "" & bh3_w7_5 & bh3_w7_6 & bh3_w7_0 & bh3_w7_1 & bh3_w7_2 & bh3_w7_3;
   bh3_w7_9 <= Compressor_6_3_comb_uid209_bh3_uid249_Out0(0);
   bh3_w8_5 <= Compressor_6_3_comb_uid209_bh3_uid249_Out0(1);
   bh3_w9_4 <= Compressor_6_3_comb_uid209_bh3_uid249_Out0(2);
   Compressor_6_3_comb_uid209_uid249: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid249_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid249_Out0);


   Compressor_14_3_comb_uid204_bh3_uid250_In0 <= "" & bh3_w8_3 & bh3_w8_0 & bh3_w8_1 & bh3_w8_2;
   Compressor_14_3_comb_uid204_bh3_uid250_In1 <= "" & bh3_w9_3;
   bh3_w8_6 <= Compressor_14_3_comb_uid204_bh3_uid250_Out0(0);
   bh3_w9_5 <= Compressor_14_3_comb_uid204_bh3_uid250_Out0(1);
   bh3_w10_3 <= Compressor_14_3_comb_uid204_bh3_uid250_Out0(2);
   Compressor_14_3_comb_uid204_uid250: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid250_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid250_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid250_Out0);


   Compressor_23_3_comb_uid198_bh3_uid251_In0 <= "" & bh3_w9_0 & bh3_w9_1 & bh3_w9_2;
   Compressor_23_3_comb_uid198_bh3_uid251_In1 <= "" & "0" & "0";
   bh3_w9_6 <= Compressor_23_3_comb_uid198_bh3_uid251_Out0(0);
   bh3_w10_4 <= Compressor_23_3_comb_uid198_bh3_uid251_Out0(1);
   bh3_w11_2 <= Compressor_23_3_comb_uid198_bh3_uid251_Out0(2);
   Compressor_23_3_comb_uid198_uid251: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid251_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid251_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid251_Out0);


   Compressor_23_3_comb_uid198_bh3_uid252_In0 <= "" & bh3_w10_2 & bh3_w10_0 & bh3_w10_1;
   Compressor_23_3_comb_uid198_bh3_uid252_In1 <= "" & bh3_w11_1 & bh3_w11_0;
   bh3_w10_5 <= Compressor_23_3_comb_uid198_bh3_uid252_Out0(0);
   bh3_w11_3 <= Compressor_23_3_comb_uid198_bh3_uid252_Out0(1);
   Compressor_23_3_comb_uid198_uid252: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid252_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid252_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid252_Out0);


   Compressor_23_3_comb_uid198_bh3_uid253_In0 <= "" & bh3_wm18_4 & bh3_wm18_3 & "0";
   Compressor_23_3_comb_uid198_bh3_uid253_In1 <= "" & bh3_wm17_5 & bh3_wm17_4;
   bh3_wm18_5 <= Compressor_23_3_comb_uid198_bh3_uid253_Out0(0);
   bh3_wm17_6 <= Compressor_23_3_comb_uid198_bh3_uid253_Out0(1);
   bh3_wm16_7 <= Compressor_23_3_comb_uid198_bh3_uid253_Out0(2);
   Compressor_23_3_comb_uid198_uid253: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid253_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid253_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid253_Out0);


   Compressor_3_2_comb_uid201_bh3_uid254_In0 <= "" & bh3_wm16_6 & bh3_wm16_5 & "0";
   bh3_wm16_8 <= Compressor_3_2_comb_uid201_bh3_uid254_Out0(0);
   bh3_wm15_8 <= Compressor_3_2_comb_uid201_bh3_uid254_Out0(1);
   Compressor_3_2_comb_uid201_uid254: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid254_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid254_Out0);


   Compressor_23_3_comb_uid198_bh3_uid255_In0 <= "" & bh3_wm15_7 & bh3_wm15_6 & bh3_wm15_5;
   Compressor_23_3_comb_uid198_bh3_uid255_In1 <= "" & bh3_wm14_8 & bh3_wm14_7;
   bh3_wm15_9 <= Compressor_23_3_comb_uid198_bh3_uid255_Out0(0);
   bh3_wm14_10 <= Compressor_23_3_comb_uid198_bh3_uid255_Out0(1);
   bh3_wm13_11 <= Compressor_23_3_comb_uid198_bh3_uid255_Out0(2);
   Compressor_23_3_comb_uid198_uid255: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid255_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid255_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid255_Out0);


   Compressor_14_3_comb_uid204_bh3_uid256_In0 <= "" & bh3_wm13_10 & bh3_wm13_7 & bh3_wm13_9 & bh3_wm13_8;
   Compressor_14_3_comb_uid204_bh3_uid256_In1 <= "" & bh3_wm12_10;
   bh3_wm13_12 <= Compressor_14_3_comb_uid204_bh3_uid256_Out0(0);
   bh3_wm12_12 <= Compressor_14_3_comb_uid204_bh3_uid256_Out0(1);
   bh3_wm11_14 <= Compressor_14_3_comb_uid204_bh3_uid256_Out0(2);
   Compressor_14_3_comb_uid204_uid256: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid256_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid256_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid256_Out0);


   Compressor_3_2_comb_uid201_bh3_uid257_In0 <= "" & bh3_wm12_11 & bh3_wm12_9 & bh3_wm12_8;
   bh3_wm12_13 <= Compressor_3_2_comb_uid201_bh3_uid257_Out0(0);
   bh3_wm11_15 <= Compressor_3_2_comb_uid201_bh3_uid257_Out0(1);
   Compressor_3_2_comb_uid201_uid257: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid257_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid257_Out0);


   Compressor_14_3_comb_uid204_bh3_uid258_In0 <= "" & bh3_wm11_13 & bh3_wm11_10 & bh3_wm11_12 & bh3_wm11_11;
   Compressor_14_3_comb_uid204_bh3_uid258_In1 <= "" & bh3_wm10_14;
   bh3_wm11_16 <= Compressor_14_3_comb_uid204_bh3_uid258_Out0(0);
   bh3_wm10_15 <= Compressor_14_3_comb_uid204_bh3_uid258_Out0(1);
   bh3_wm9_15 <= Compressor_14_3_comb_uid204_bh3_uid258_Out0(2);
   Compressor_14_3_comb_uid204_uid258: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid258_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid258_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid258_Out0);


   Compressor_14_3_comb_uid204_bh3_uid259_In0 <= "" & bh3_wm10_12 & bh3_wm10_13 & bh3_wm10_11 & bh3_wm10_10;
   Compressor_14_3_comb_uid204_bh3_uid259_In1 <= "" & bh3_wm9_14;
   bh3_wm10_16 <= Compressor_14_3_comb_uid204_bh3_uid259_Out0(0);
   bh3_wm9_16 <= Compressor_14_3_comb_uid204_bh3_uid259_Out0(1);
   bh3_wm8_18 <= Compressor_14_3_comb_uid204_bh3_uid259_Out0(2);
   Compressor_14_3_comb_uid204_uid259: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid259_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid259_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid259_Out0);


   Compressor_3_2_comb_uid201_bh3_uid260_In0 <= "" & bh3_wm9_12 & bh3_wm9_13 & bh3_wm9_11;
   bh3_wm9_17 <= Compressor_3_2_comb_uid201_bh3_uid260_Out0(0);
   bh3_wm8_19 <= Compressor_3_2_comb_uid201_bh3_uid260_Out0(1);
   Compressor_3_2_comb_uid201_uid260: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid260_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid260_Out0);


   Compressor_6_3_comb_uid209_bh3_uid261_In0 <= "" & bh3_wm8_15 & bh3_wm8_13 & bh3_wm8_16 & bh3_wm8_14 & bh3_wm8_12 & bh3_wm8_17;
   bh3_wm8_20 <= Compressor_6_3_comb_uid209_bh3_uid261_Out0(0);
   bh3_wm7_17 <= Compressor_6_3_comb_uid209_bh3_uid261_Out0(1);
   bh3_wm6_19 <= Compressor_6_3_comb_uid209_bh3_uid261_Out0(2);
   Compressor_6_3_comb_uid209_uid261: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid261_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid261_Out0);


   Compressor_14_3_comb_uid204_bh3_uid262_In0 <= "" & bh3_wm7_12 & bh3_wm7_13 & bh3_wm7_14 & bh3_wm7_15;
   Compressor_14_3_comb_uid204_bh3_uid262_In1 <= "" & bh3_wm6_11;
   bh3_wm7_18 <= Compressor_14_3_comb_uid204_bh3_uid262_Out0(0);
   bh3_wm6_20 <= Compressor_14_3_comb_uid204_bh3_uid262_Out0(1);
   bh3_wm5_21 <= Compressor_14_3_comb_uid204_bh3_uid262_Out0(2);
   Compressor_14_3_comb_uid204_uid262: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid262_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid262_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid262_Out0);


   Compressor_6_3_comb_uid209_bh3_uid263_In0 <= "" & bh3_wm6_17 & bh3_wm6_13 & bh3_wm6_14 & bh3_wm6_15 & bh3_wm6_16 & bh3_wm6_18;
   bh3_wm6_21 <= Compressor_6_3_comb_uid209_bh3_uid263_Out0(0);
   bh3_wm5_22 <= Compressor_6_3_comb_uid209_bh3_uid263_Out0(1);
   bh3_wm4_21 <= Compressor_6_3_comb_uid209_bh3_uid263_Out0(2);
   Compressor_6_3_comb_uid209_uid263: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid263_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid263_Out0);


   Compressor_6_3_comb_uid209_bh3_uid264_In0 <= "" & bh3_wm5_20 & bh3_wm5_18 & bh3_wm5_16 & bh3_wm5_15 & bh3_wm5_14 & bh3_wm5_17;
   bh3_wm5_23 <= Compressor_6_3_comb_uid209_bh3_uid264_Out0(0);
   bh3_wm4_22 <= Compressor_6_3_comb_uid209_bh3_uid264_Out0(1);
   bh3_wm3_23 <= Compressor_6_3_comb_uid209_bh3_uid264_Out0(2);
   Compressor_6_3_comb_uid209_uid264: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid264_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid264_Out0);


   Compressor_6_3_comb_uid209_bh3_uid265_In0 <= "" & bh3_wm4_18 & bh3_wm4_19 & bh3_wm4_16 & bh3_wm4_15 & bh3_wm4_14 & bh3_wm4_17;
   bh3_wm4_23 <= Compressor_6_3_comb_uid209_bh3_uid265_Out0(0);
   bh3_wm3_24 <= Compressor_6_3_comb_uid209_bh3_uid265_Out0(1);
   bh3_wm2_20 <= Compressor_6_3_comb_uid209_bh3_uid265_Out0(2);
   Compressor_6_3_comb_uid209_uid265: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid265_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid265_Out0);


   Compressor_6_3_comb_uid209_bh3_uid266_In0 <= "" & bh3_wm3_22 & bh3_wm3_17 & bh3_wm3_21 & bh3_wm3_20 & bh3_wm3_19 & "0";
   bh3_wm3_25 <= Compressor_6_3_comb_uid209_bh3_uid266_Out0(0);
   bh3_wm2_21 <= Compressor_6_3_comb_uid209_bh3_uid266_Out0(1);
   bh3_wm1_18 <= Compressor_6_3_comb_uid209_bh3_uid266_Out0(2);
   Compressor_6_3_comb_uid209_uid266: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid266_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid266_Out0);


   Compressor_23_3_comb_uid198_bh3_uid267_In0 <= "" & bh3_wm3_18 & bh3_wm3_16 & bh3_wm3_15;
   Compressor_23_3_comb_uid198_bh3_uid267_In1 <= "" & bh3_wm2_11 & bh3_wm2_17;
   bh3_wm3_26 <= Compressor_23_3_comb_uid198_bh3_uid267_Out0(0);
   bh3_wm2_22 <= Compressor_23_3_comb_uid198_bh3_uid267_Out0(1);
   bh3_wm1_19 <= Compressor_23_3_comb_uid198_bh3_uid267_Out0(2);
   Compressor_23_3_comb_uid198_uid267: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid267_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid267_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid267_Out0);


   Compressor_6_3_comb_uid209_bh3_uid268_In0 <= "" & bh3_wm2_18 & bh3_wm2_13 & bh3_wm2_14 & bh3_wm2_15 & bh3_wm2_16 & bh3_wm2_19;
   bh3_wm2_23 <= Compressor_6_3_comb_uid209_bh3_uid268_Out0(0);
   bh3_wm1_20 <= Compressor_6_3_comb_uid209_bh3_uid268_Out0(1);
   bh3_w0_18 <= Compressor_6_3_comb_uid209_bh3_uid268_Out0(2);
   Compressor_6_3_comb_uid209_uid268: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid268_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid268_Out0);


   Compressor_6_3_comb_uid209_bh3_uid269_In0 <= "" & bh3_wm1_16 & bh3_wm1_15 & bh3_wm1_14 & bh3_wm1_13 & bh3_wm1_12 & bh3_wm1_17;
   bh3_wm1_21 <= Compressor_6_3_comb_uid209_bh3_uid269_Out0(0);
   bh3_w0_19 <= Compressor_6_3_comb_uid209_bh3_uid269_Out0(1);
   bh3_w1_18 <= Compressor_6_3_comb_uid209_bh3_uid269_Out0(2);
   Compressor_6_3_comb_uid209_uid269: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid269_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid269_Out0);


   Compressor_6_3_comb_uid209_bh3_uid270_In0 <= "" & bh3_w0_17 & bh3_w0_16 & bh3_w0_15 & bh3_w0_14 & bh3_w0_13 & bh3_w0_12;
   bh3_w0_20 <= Compressor_6_3_comb_uid209_bh3_uid270_Out0(0);
   bh3_w1_19 <= Compressor_6_3_comb_uid209_bh3_uid270_Out0(1);
   bh3_w2_15 <= Compressor_6_3_comb_uid209_bh3_uid270_Out0(2);
   Compressor_6_3_comb_uid209_uid270: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid270_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid270_Out0);


   Compressor_6_3_comb_uid209_bh3_uid271_In0 <= "" & bh3_w1_17 & bh3_w1_16 & bh3_w1_15 & bh3_w1_14 & bh3_w1_13 & bh3_w1_12;
   bh3_w1_20 <= Compressor_6_3_comb_uid209_bh3_uid271_Out0(0);
   bh3_w2_16 <= Compressor_6_3_comb_uid209_bh3_uid271_Out0(1);
   bh3_w3_14 <= Compressor_6_3_comb_uid209_bh3_uid271_Out0(2);
   Compressor_6_3_comb_uid209_uid271: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid271_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid271_Out0);


   Compressor_6_3_comb_uid209_bh3_uid272_In0 <= "" & bh3_w2_14 & bh3_w2_13 & bh3_w2_12 & bh3_w2_11 & bh3_w2_10 & bh3_w2_9;
   bh3_w2_17 <= Compressor_6_3_comb_uid209_bh3_uid272_Out0(0);
   bh3_w3_15 <= Compressor_6_3_comb_uid209_bh3_uid272_Out0(1);
   bh3_w4_13 <= Compressor_6_3_comb_uid209_bh3_uid272_Out0(2);
   Compressor_6_3_comb_uid209_uid272: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid272_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid272_Out0);


   Compressor_6_3_comb_uid209_bh3_uid273_In0 <= "" & bh3_w3_7 & bh3_w3_12 & bh3_w3_13 & bh3_w3_11 & bh3_w3_10 & bh3_w3_9;
   bh3_w3_16 <= Compressor_6_3_comb_uid209_bh3_uid273_Out0(0);
   bh3_w4_14 <= Compressor_6_3_comb_uid209_bh3_uid273_Out0(1);
   bh3_w5_11 <= Compressor_6_3_comb_uid209_bh3_uid273_Out0(2);
   Compressor_6_3_comb_uid209_uid273: Compressor_6_3_comb_uid209
      port map ( X0 => Compressor_6_3_comb_uid209_bh3_uid273_In0,
                 R => Compressor_6_3_comb_uid209_bh3_uid273_Out0);


   Compressor_14_3_comb_uid204_bh3_uid274_In0 <= "" & bh3_w4_12 & bh3_w4_9 & bh3_w4_11 & bh3_w4_10;
   Compressor_14_3_comb_uid204_bh3_uid274_In1 <= "" & bh3_w5_9;
   bh3_w4_15 <= Compressor_14_3_comb_uid204_bh3_uid274_Out0(0);
   bh3_w5_12 <= Compressor_14_3_comb_uid204_bh3_uid274_Out0(1);
   bh3_w6_11 <= Compressor_14_3_comb_uid204_bh3_uid274_Out0(2);
   Compressor_14_3_comb_uid204_uid274: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid274_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid274_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid274_Out0);


   Compressor_3_2_comb_uid201_bh3_uid275_In0 <= "" & bh3_w5_10 & bh3_w5_8 & bh3_w5_7;
   bh3_w5_13 <= Compressor_3_2_comb_uid201_bh3_uid275_Out0(0);
   bh3_w6_12 <= Compressor_3_2_comb_uid201_bh3_uid275_Out0(1);
   Compressor_3_2_comb_uid201_uid275: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid275_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid275_Out0);


   Compressor_14_3_comb_uid204_bh3_uid276_In0 <= "" & bh3_w6_4 & bh3_w6_8 & bh3_w6_10 & bh3_w6_9;
   Compressor_14_3_comb_uid204_bh3_uid276_In1 <= "" & bh3_w7_4;
   bh3_w6_13 <= Compressor_14_3_comb_uid204_bh3_uid276_Out0(0);
   bh3_w7_10 <= Compressor_14_3_comb_uid204_bh3_uid276_Out0(1);
   bh3_w8_7 <= Compressor_14_3_comb_uid204_bh3_uid276_Out0(2);
   Compressor_14_3_comb_uid204_uid276: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid276_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid276_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid276_Out0);


   Compressor_23_3_comb_uid198_bh3_uid277_In0 <= "" & bh3_w7_9 & bh3_w7_8 & bh3_w7_7;
   Compressor_23_3_comb_uid198_bh3_uid277_In1 <= "" & bh3_w8_6 & bh3_w8_5;
   bh3_w7_11 <= Compressor_23_3_comb_uid198_bh3_uid277_Out0(0);
   bh3_w8_8 <= Compressor_23_3_comb_uid198_bh3_uid277_Out0(1);
   bh3_w9_7 <= Compressor_23_3_comb_uid198_bh3_uid277_Out0(2);
   Compressor_23_3_comb_uid198_uid277: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid277_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid277_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid277_Out0);


   Compressor_23_3_comb_uid198_bh3_uid278_In0 <= "" & bh3_w9_6 & bh3_w9_5 & bh3_w9_4;
   Compressor_23_3_comb_uid198_bh3_uid278_In1 <= "" & bh3_w10_5 & bh3_w10_4;
   bh3_w9_8 <= Compressor_23_3_comb_uid198_bh3_uid278_Out0(0);
   bh3_w10_6 <= Compressor_23_3_comb_uid198_bh3_uid278_Out0(1);
   bh3_w11_4 <= Compressor_23_3_comb_uid198_bh3_uid278_Out0(2);
   Compressor_23_3_comb_uid198_uid278: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid278_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid278_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid278_Out0);


   Compressor_14_3_comb_uid204_bh3_uid279_In0 <= "" & bh3_w11_3 & bh3_w11_2 & "0" & "0";
   Compressor_14_3_comb_uid204_bh3_uid279_In1 <= "" & "0";
   bh3_w11_5 <= Compressor_14_3_comb_uid204_bh3_uid279_Out0(0);
   Compressor_14_3_comb_uid204_uid279: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid279_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid279_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid279_Out0);


   Compressor_23_3_comb_uid198_bh3_uid280_In0 <= "" & bh3_wm16_8 & bh3_wm16_7 & "0";
   Compressor_23_3_comb_uid198_bh3_uid280_In1 <= "" & bh3_wm15_9 & bh3_wm15_8;
   bh3_wm16_9 <= Compressor_23_3_comb_uid198_bh3_uid280_Out0(0);
   bh3_wm15_10 <= Compressor_23_3_comb_uid198_bh3_uid280_Out0(1);
   bh3_wm14_11 <= Compressor_23_3_comb_uid198_bh3_uid280_Out0(2);
   Compressor_23_3_comb_uid198_uid280: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid280_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid280_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid280_Out0);


   Compressor_23_3_comb_uid198_bh3_uid281_In0 <= "" & bh3_wm14_9 & bh3_wm14_10 & "0";
   Compressor_23_3_comb_uid198_bh3_uid281_In1 <= "" & bh3_wm13_11 & bh3_wm13_12;
   bh3_wm14_12 <= Compressor_23_3_comb_uid198_bh3_uid281_Out0(0);
   bh3_wm13_13 <= Compressor_23_3_comb_uid198_bh3_uid281_Out0(1);
   bh3_wm12_14 <= Compressor_23_3_comb_uid198_bh3_uid281_Out0(2);
   Compressor_23_3_comb_uid198_uid281: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid281_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid281_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid281_Out0);


   Compressor_3_2_comb_uid201_bh3_uid282_In0 <= "" & bh3_wm12_13 & bh3_wm12_12 & "0";
   bh3_wm12_15 <= Compressor_3_2_comb_uid201_bh3_uid282_Out0(0);
   bh3_wm11_17 <= Compressor_3_2_comb_uid201_bh3_uid282_Out0(1);
   Compressor_3_2_comb_uid201_uid282: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid282_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid282_Out0);


   Compressor_14_3_comb_uid204_bh3_uid283_In0 <= "" & bh3_wm11_9 & bh3_wm11_16 & bh3_wm11_15 & bh3_wm11_14;
   Compressor_14_3_comb_uid204_bh3_uid283_In1 <= "" & bh3_wm10_16;
   bh3_wm11_18 <= Compressor_14_3_comb_uid204_bh3_uid283_Out0(0);
   bh3_wm10_17 <= Compressor_14_3_comb_uid204_bh3_uid283_Out0(1);
   bh3_wm9_18 <= Compressor_14_3_comb_uid204_bh3_uid283_Out0(2);
   Compressor_14_3_comb_uid204_uid283: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid283_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid283_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid283_Out0);


   Compressor_14_3_comb_uid204_bh3_uid284_In0 <= "" & bh3_wm9_10 & bh3_wm9_17 & bh3_wm9_16 & bh3_wm9_15;
   Compressor_14_3_comb_uid204_bh3_uid284_In1 <= "" & "0";
   bh3_wm9_19 <= Compressor_14_3_comb_uid204_bh3_uid284_Out0(0);
   bh3_wm8_21 <= Compressor_14_3_comb_uid204_bh3_uid284_Out0(1);
   bh3_wm7_19 <= Compressor_14_3_comb_uid204_bh3_uid284_Out0(2);
   Compressor_14_3_comb_uid204_uid284: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid284_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid284_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid284_Out0);


   Compressor_3_2_comb_uid201_bh3_uid285_In0 <= "" & bh3_wm8_19 & bh3_wm8_18 & bh3_wm8_20;
   bh3_wm8_22 <= Compressor_3_2_comb_uid201_bh3_uid285_Out0(0);
   bh3_wm7_20 <= Compressor_3_2_comb_uid201_bh3_uid285_Out0(1);
   Compressor_3_2_comb_uid201_uid285: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid285_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid285_Out0);


   Compressor_23_3_comb_uid198_bh3_uid286_In0 <= "" & bh3_wm7_16 & bh3_wm7_18 & bh3_wm7_17;
   Compressor_23_3_comb_uid198_bh3_uid286_In1 <= "" & bh3_wm6_20 & bh3_wm6_21;
   bh3_wm7_21 <= Compressor_23_3_comb_uid198_bh3_uid286_Out0(0);
   bh3_wm6_22 <= Compressor_23_3_comb_uid198_bh3_uid286_Out0(1);
   bh3_wm5_24 <= Compressor_23_3_comb_uid198_bh3_uid286_Out0(2);
   Compressor_23_3_comb_uid198_uid286: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid286_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid286_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid286_Out0);


   Compressor_14_3_comb_uid204_bh3_uid287_In0 <= "" & bh3_wm5_19 & bh3_wm5_21 & bh3_wm5_23 & bh3_wm5_22;
   Compressor_14_3_comb_uid204_bh3_uid287_In1 <= "" & bh3_wm4_20;
   bh3_wm5_25 <= Compressor_14_3_comb_uid204_bh3_uid287_Out0(0);
   bh3_wm4_24 <= Compressor_14_3_comb_uid204_bh3_uid287_Out0(1);
   bh3_wm3_27 <= Compressor_14_3_comb_uid204_bh3_uid287_Out0(2);
   Compressor_14_3_comb_uid204_uid287: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid287_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid287_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid287_Out0);


   Compressor_3_2_comb_uid201_bh3_uid288_In0 <= "" & bh3_wm4_23 & bh3_wm4_22 & bh3_wm4_21;
   bh3_wm4_25 <= Compressor_3_2_comb_uid201_bh3_uid288_Out0(0);
   bh3_wm3_28 <= Compressor_3_2_comb_uid201_bh3_uid288_Out0(1);
   Compressor_3_2_comb_uid201_uid288: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid288_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid288_Out0);


   Compressor_14_3_comb_uid204_bh3_uid289_In0 <= "" & bh3_wm3_26 & bh3_wm3_25 & bh3_wm3_24 & bh3_wm3_23;
   Compressor_14_3_comb_uid204_bh3_uid289_In1 <= "" & bh3_wm2_22;
   bh3_wm3_29 <= Compressor_14_3_comb_uid204_bh3_uid289_Out0(0);
   bh3_wm2_24 <= Compressor_14_3_comb_uid204_bh3_uid289_Out0(1);
   bh3_wm1_22 <= Compressor_14_3_comb_uid204_bh3_uid289_Out0(2);
   Compressor_14_3_comb_uid204_uid289: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid289_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid289_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid289_Out0);


   Compressor_3_2_comb_uid201_bh3_uid290_In0 <= "" & bh3_wm2_23 & bh3_wm2_21 & bh3_wm2_20;
   bh3_wm2_25 <= Compressor_3_2_comb_uid201_bh3_uid290_Out0(0);
   bh3_wm1_23 <= Compressor_3_2_comb_uid201_bh3_uid290_Out0(1);
   Compressor_3_2_comb_uid201_uid290: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid290_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid290_Out0);


   Compressor_14_3_comb_uid204_bh3_uid291_In0 <= "" & bh3_wm1_19 & bh3_wm1_21 & bh3_wm1_20 & bh3_wm1_18;
   Compressor_14_3_comb_uid204_bh3_uid291_In1 <= "" & "0";
   bh3_wm1_24 <= Compressor_14_3_comb_uid204_bh3_uid291_Out0(0);
   bh3_w0_21 <= Compressor_14_3_comb_uid204_bh3_uid291_Out0(1);
   bh3_w1_21 <= Compressor_14_3_comb_uid204_bh3_uid291_Out0(2);
   Compressor_14_3_comb_uid204_uid291: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid291_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid291_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid291_Out0);


   Compressor_3_2_comb_uid201_bh3_uid292_In0 <= "" & bh3_w0_20 & bh3_w0_19 & bh3_w0_18;
   bh3_w0_22 <= Compressor_3_2_comb_uid201_bh3_uid292_Out0(0);
   bh3_w1_22 <= Compressor_3_2_comb_uid201_bh3_uid292_Out0(1);
   Compressor_3_2_comb_uid201_uid292: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid292_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid292_Out0);


   Compressor_23_3_comb_uid198_bh3_uid293_In0 <= "" & bh3_w1_20 & bh3_w1_19 & bh3_w1_18;
   Compressor_23_3_comb_uid198_bh3_uid293_In1 <= "" & bh3_w2_17 & bh3_w2_16;
   bh3_w1_23 <= Compressor_23_3_comb_uid198_bh3_uid293_Out0(0);
   bh3_w2_18 <= Compressor_23_3_comb_uid198_bh3_uid293_Out0(1);
   bh3_w3_17 <= Compressor_23_3_comb_uid198_bh3_uid293_Out0(2);
   Compressor_23_3_comb_uid198_uid293: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid293_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid293_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid293_Out0);


   Compressor_3_2_comb_uid201_bh3_uid294_In0 <= "" & bh3_w3_16 & bh3_w3_15 & bh3_w3_14;
   bh3_w3_18 <= Compressor_3_2_comb_uid201_bh3_uid294_Out0(0);
   bh3_w4_16 <= Compressor_3_2_comb_uid201_bh3_uid294_Out0(1);
   Compressor_3_2_comb_uid201_uid294: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid294_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid294_Out0);


   Compressor_14_3_comb_uid204_bh3_uid295_In0 <= "" & bh3_w4_8 & bh3_w4_15 & bh3_w4_14 & bh3_w4_13;
   Compressor_14_3_comb_uid204_bh3_uid295_In1 <= "" & "0";
   bh3_w4_17 <= Compressor_14_3_comb_uid204_bh3_uid295_Out0(0);
   bh3_w5_14 <= Compressor_14_3_comb_uid204_bh3_uid295_Out0(1);
   bh3_w6_14 <= Compressor_14_3_comb_uid204_bh3_uid295_Out0(2);
   Compressor_14_3_comb_uid204_uid295: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid295_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid295_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid295_Out0);


   Compressor_3_2_comb_uid201_bh3_uid296_In0 <= "" & bh3_w5_13 & bh3_w5_12 & bh3_w5_11;
   bh3_w5_15 <= Compressor_3_2_comb_uid201_bh3_uid296_Out0(0);
   bh3_w6_15 <= Compressor_3_2_comb_uid201_bh3_uid296_Out0(1);
   Compressor_3_2_comb_uid201_uid296: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid296_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid296_Out0);


   Compressor_14_3_comb_uid204_bh3_uid297_In0 <= "" & bh3_w6_7 & bh3_w6_13 & bh3_w6_12 & bh3_w6_11;
   Compressor_14_3_comb_uid204_bh3_uid297_In1 <= "" & bh3_w7_11;
   bh3_w6_16 <= Compressor_14_3_comb_uid204_bh3_uid297_Out0(0);
   bh3_w7_12 <= Compressor_14_3_comb_uid204_bh3_uid297_Out0(1);
   bh3_w8_9 <= Compressor_14_3_comb_uid204_bh3_uid297_Out0(2);
   Compressor_14_3_comb_uid204_uid297: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid297_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid297_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid297_Out0);


   Compressor_23_3_comb_uid198_bh3_uid298_In0 <= "" & bh3_w8_4 & bh3_w8_8 & bh3_w8_7;
   Compressor_23_3_comb_uid198_bh3_uid298_In1 <= "" & bh3_w9_8 & bh3_w9_7;
   bh3_w8_10 <= Compressor_23_3_comb_uid198_bh3_uid298_Out0(0);
   bh3_w9_9 <= Compressor_23_3_comb_uid198_bh3_uid298_Out0(1);
   bh3_w10_7 <= Compressor_23_3_comb_uid198_bh3_uid298_Out0(2);
   Compressor_23_3_comb_uid198_uid298: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid298_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid298_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid298_Out0);


   Compressor_23_3_comb_uid198_bh3_uid299_In0 <= "" & bh3_w10_3 & bh3_w10_6 & "0";
   Compressor_23_3_comb_uid198_bh3_uid299_In1 <= "" & bh3_w11_5 & bh3_w11_4;
   bh3_w10_8 <= Compressor_23_3_comb_uid198_bh3_uid299_Out0(0);
   bh3_w11_6 <= Compressor_23_3_comb_uid198_bh3_uid299_Out0(1);
   Compressor_23_3_comb_uid198_uid299: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid299_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid299_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid299_Out0);


   Compressor_14_3_comb_uid204_bh3_uid300_In0 <= "" & bh3_wm14_11 & bh3_wm14_12 & "0" & "0";
   Compressor_14_3_comb_uid204_bh3_uid300_In1 <= "" & bh3_wm13_13;
   bh3_wm14_13 <= Compressor_14_3_comb_uid204_bh3_uid300_Out0(0);
   bh3_wm13_14 <= Compressor_14_3_comb_uid204_bh3_uid300_Out0(1);
   bh3_wm12_16 <= Compressor_14_3_comb_uid204_bh3_uid300_Out0(2);
   Compressor_14_3_comb_uid204_uid300: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid300_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid300_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid300_Out0);


   Compressor_23_3_comb_uid198_bh3_uid301_In0 <= "" & bh3_wm12_15 & bh3_wm12_14 & "0";
   Compressor_23_3_comb_uid198_bh3_uid301_In1 <= "" & bh3_wm11_18 & bh3_wm11_17;
   bh3_wm12_17 <= Compressor_23_3_comb_uid198_bh3_uid301_Out0(0);
   bh3_wm11_19 <= Compressor_23_3_comb_uid198_bh3_uid301_Out0(1);
   bh3_wm10_18 <= Compressor_23_3_comb_uid198_bh3_uid301_Out0(2);
   Compressor_23_3_comb_uid198_uid301: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid301_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid301_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid301_Out0);


   Compressor_23_3_comb_uid198_bh3_uid302_In0 <= "" & bh3_wm10_15 & bh3_wm10_17 & "0";
   Compressor_23_3_comb_uid198_bh3_uid302_In1 <= "" & bh3_wm9_19 & bh3_wm9_18;
   bh3_wm10_19 <= Compressor_23_3_comb_uid198_bh3_uid302_Out0(0);
   bh3_wm9_20 <= Compressor_23_3_comb_uid198_bh3_uid302_Out0(1);
   bh3_wm8_23 <= Compressor_23_3_comb_uid198_bh3_uid302_Out0(2);
   Compressor_23_3_comb_uid198_uid302: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid302_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid302_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid302_Out0);


   Compressor_3_2_comb_uid201_bh3_uid303_In0 <= "" & bh3_wm8_21 & bh3_wm8_22 & "0";
   bh3_wm8_24 <= Compressor_3_2_comb_uid201_bh3_uid303_Out0(0);
   bh3_wm7_22 <= Compressor_3_2_comb_uid201_bh3_uid303_Out0(1);
   Compressor_3_2_comb_uid201_uid303: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid303_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid303_Out0);


   Compressor_23_3_comb_uid198_bh3_uid304_In0 <= "" & bh3_wm7_19 & bh3_wm7_21 & bh3_wm7_20;
   Compressor_23_3_comb_uid198_bh3_uid304_In1 <= "" & bh3_wm6_19 & bh3_wm6_22;
   bh3_wm7_23 <= Compressor_23_3_comb_uid198_bh3_uid304_Out0(0);
   bh3_wm6_23 <= Compressor_23_3_comb_uid198_bh3_uid304_Out0(1);
   bh3_wm5_26 <= Compressor_23_3_comb_uid198_bh3_uid304_Out0(2);
   Compressor_23_3_comb_uid198_uid304: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid304_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid304_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid304_Out0);


   Compressor_23_3_comb_uid198_bh3_uid305_In0 <= "" & bh3_wm5_25 & bh3_wm5_24 & "0";
   Compressor_23_3_comb_uid198_bh3_uid305_In1 <= "" & bh3_wm4_25 & bh3_wm4_24;
   bh3_wm5_27 <= Compressor_23_3_comb_uid198_bh3_uid305_Out0(0);
   bh3_wm4_26 <= Compressor_23_3_comb_uid198_bh3_uid305_Out0(1);
   bh3_wm3_30 <= Compressor_23_3_comb_uid198_bh3_uid305_Out0(2);
   Compressor_23_3_comb_uid198_uid305: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid305_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid305_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid305_Out0);


   Compressor_23_3_comb_uid198_bh3_uid306_In0 <= "" & bh3_wm3_29 & bh3_wm3_28 & bh3_wm3_27;
   Compressor_23_3_comb_uid198_bh3_uid306_In1 <= "" & bh3_wm2_25 & bh3_wm2_24;
   bh3_wm3_31 <= Compressor_23_3_comb_uid198_bh3_uid306_Out0(0);
   bh3_wm2_26 <= Compressor_23_3_comb_uid198_bh3_uid306_Out0(1);
   bh3_wm1_25 <= Compressor_23_3_comb_uid198_bh3_uid306_Out0(2);
   Compressor_23_3_comb_uid198_uid306: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid306_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid306_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid306_Out0);


   Compressor_23_3_comb_uid198_bh3_uid307_In0 <= "" & bh3_wm1_24 & bh3_wm1_23 & bh3_wm1_22;
   Compressor_23_3_comb_uid198_bh3_uid307_In1 <= "" & bh3_w0_22 & bh3_w0_21;
   bh3_wm1_26 <= Compressor_23_3_comb_uid198_bh3_uid307_Out0(0);
   bh3_w0_23 <= Compressor_23_3_comb_uid198_bh3_uid307_Out0(1);
   bh3_w1_24 <= Compressor_23_3_comb_uid198_bh3_uid307_Out0(2);
   Compressor_23_3_comb_uid198_uid307: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid307_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid307_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid307_Out0);


   Compressor_23_3_comb_uid198_bh3_uid308_In0 <= "" & bh3_w1_23 & bh3_w1_22 & bh3_w1_21;
   Compressor_23_3_comb_uid198_bh3_uid308_In1 <= "" & bh3_w2_15 & bh3_w2_18;
   bh3_w1_25 <= Compressor_23_3_comb_uid198_bh3_uid308_Out0(0);
   bh3_w2_19 <= Compressor_23_3_comb_uid198_bh3_uid308_Out0(1);
   bh3_w3_19 <= Compressor_23_3_comb_uid198_bh3_uid308_Out0(2);
   Compressor_23_3_comb_uid198_uid308: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid308_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid308_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid308_Out0);


   Compressor_23_3_comb_uid198_bh3_uid309_In0 <= "" & bh3_w3_18 & bh3_w3_17 & "0";
   Compressor_23_3_comb_uid198_bh3_uid309_In1 <= "" & bh3_w4_17 & bh3_w4_16;
   bh3_w3_20 <= Compressor_23_3_comb_uid198_bh3_uid309_Out0(0);
   bh3_w4_18 <= Compressor_23_3_comb_uid198_bh3_uid309_Out0(1);
   bh3_w5_16 <= Compressor_23_3_comb_uid198_bh3_uid309_Out0(2);
   Compressor_23_3_comb_uid198_uid309: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid309_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid309_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid309_Out0);


   Compressor_3_2_comb_uid201_bh3_uid310_In0 <= "" & bh3_w5_15 & bh3_w5_14 & "0";
   bh3_w5_17 <= Compressor_3_2_comb_uid201_bh3_uid310_Out0(0);
   bh3_w6_17 <= Compressor_3_2_comb_uid201_bh3_uid310_Out0(1);
   Compressor_3_2_comb_uid201_uid310: Compressor_3_2_comb_uid201
      port map ( X0 => Compressor_3_2_comb_uid201_bh3_uid310_In0,
                 R => Compressor_3_2_comb_uid201_bh3_uid310_Out0);


   Compressor_23_3_comb_uid198_bh3_uid311_In0 <= "" & bh3_w6_16 & bh3_w6_15 & bh3_w6_14;
   Compressor_23_3_comb_uid198_bh3_uid311_In1 <= "" & bh3_w7_10 & bh3_w7_12;
   bh3_w6_18 <= Compressor_23_3_comb_uid198_bh3_uid311_Out0(0);
   bh3_w7_13 <= Compressor_23_3_comb_uid198_bh3_uid311_Out0(1);
   bh3_w8_11 <= Compressor_23_3_comb_uid198_bh3_uid311_Out0(2);
   Compressor_23_3_comb_uid198_uid311: Compressor_23_3_comb_uid198
      port map ( X0 => Compressor_23_3_comb_uid198_bh3_uid311_In0,
                 X1 => Compressor_23_3_comb_uid198_bh3_uid311_In1,
                 R => Compressor_23_3_comb_uid198_bh3_uid311_Out0);


   Compressor_14_3_comb_uid204_bh3_uid312_In0 <= "" & bh3_w8_10 & bh3_w8_9 & "0" & "0";
   Compressor_14_3_comb_uid204_bh3_uid312_In1 <= "" & bh3_w9_9;
   bh3_w8_12 <= Compressor_14_3_comb_uid204_bh3_uid312_Out0(0);
   bh3_w9_10 <= Compressor_14_3_comb_uid204_bh3_uid312_Out0(1);
   bh3_w10_9 <= Compressor_14_3_comb_uid204_bh3_uid312_Out0(2);
   Compressor_14_3_comb_uid204_uid312: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid312_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid312_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid312_Out0);


   Compressor_14_3_comb_uid204_bh3_uid313_In0 <= "" & bh3_w10_8 & bh3_w10_7 & "0" & "0";
   Compressor_14_3_comb_uid204_bh3_uid313_In1 <= "" & bh3_w11_6;
   bh3_w10_10 <= Compressor_14_3_comb_uid204_bh3_uid313_Out0(0);
   bh3_w11_7 <= Compressor_14_3_comb_uid204_bh3_uid313_Out0(1);
   Compressor_14_3_comb_uid204_uid313: Compressor_14_3_comb_uid204
      port map ( X0 => Compressor_14_3_comb_uid204_bh3_uid313_In0,
                 X1 => Compressor_14_3_comb_uid204_bh3_uid313_In1,
                 R => Compressor_14_3_comb_uid204_bh3_uid313_Out0);

   tmp_bitheapResult_bh3_7 <= bh3_wm13_14 & bh3_wm14_13 & bh3_wm15_10 & bh3_wm16_9 & bh3_wm17_6 & bh3_wm18_5 & bh3_wm19_2 & bh3_wm20_2;

   bitheapFinalAdd_bh3_In0 <= "0" & bh3_w11_7 & bh3_w10_10 & bh3_w9_10 & bh3_w8_12 & bh3_w7_13 & bh3_w6_18 & bh3_w5_17 & bh3_w4_18 & bh3_w3_20 & bh3_w2_19 & bh3_w1_25 & bh3_w0_23 & bh3_wm1_26 & bh3_wm2_26 & bh3_wm3_31 & bh3_wm4_26 & bh3_wm5_27 & bh3_wm6_23 & bh3_wm7_23 & bh3_wm8_23 & bh3_wm9_20 & bh3_wm10_19 & bh3_wm11_19 & bh3_wm12_17;
   bitheapFinalAdd_bh3_In1 <= "0" & "0" & bh3_w10_9 & "0" & bh3_w8_11 & "0" & bh3_w6_17 & bh3_w5_16 & "0" & bh3_w3_19 & "0" & bh3_w1_24 & "0" & bh3_wm1_25 & "0" & bh3_wm3_30 & "0" & bh3_wm5_26 & "0" & bh3_wm7_22 & bh3_wm8_24 & "0" & bh3_wm10_18 & "0" & bh3_wm12_16;
   bitheapFinalAdd_bh3_Cin <= '0';

   bitheapFinalAdd_bh3: IntAdder_25_comb_uid315
      port map ( Cin => bitheapFinalAdd_bh3_Cin,
                 X => bitheapFinalAdd_bh3_In0,
                 Y => bitheapFinalAdd_bh3_In1,
                 R => bitheapFinalAdd_bh3_Out);
   bitheapResult_bh3 <= bitheapFinalAdd_bh3_Out(23 downto 0) & tmp_bitheapResult_bh3_7;
   RR <= signed(bitheapResult_bh3(31 downto 0));
R <= std_logic_vector(RR);  
end architecture;

